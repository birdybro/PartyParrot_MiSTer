/********************************************************
 * Title    : Image ROM
 * Date     : 2020/05/13
 * Design   : kingyo
 ********************************************************/
// MIT License
//
// Copyright (c) 2020 kingyo
//
// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be included in all
// copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

module ImgROM (
    input   wire            i_clk,
    input   wire            i_res_n,
    input   wire    [12:0]  i_addr,
    output  reg     [ 7:0]  o_data
    );
    
    always @(posedge i_clk or negedge i_res_n) begin
        if (~i_res_n) begin
            o_data <= 8'd0;
        end else begin
            o_data <= imageROM( i_addr );
        end
    end
    
    function [7:0] imageROM;
        input   [12:0]   addr;
        begin
            case (addr)
            // r01.bmp
                0: imageROM = 8'd63;
                1: imageROM = 8'd63;
                2: imageROM = 8'd63;
                3: imageROM = 8'd63;
                4: imageROM = 8'd63;
                5: imageROM = 8'd63;
                6: imageROM = 8'd63;
                7: imageROM = 8'd63;
                8: imageROM = 8'd63;
                9: imageROM = 8'd63;
                10: imageROM = 8'd63;
                11: imageROM = 8'd63;
                12: imageROM = 8'd63;
                13: imageROM = 8'd63;
                14: imageROM = 8'd63;
                15: imageROM = 8'd25;
                16: imageROM = 8'd77;
                17: imageROM = 8'd63;
                18: imageROM = 8'd47;
                19: imageROM = 8'd88;
                20: imageROM = 8'd63;
                21: imageROM = 8'd38;
                22: imageROM = 8'd94;
                23: imageROM = 8'd63;
                24: imageROM = 8'd33;
                25: imageROM = 8'd98;
                26: imageROM = 8'd63;
                27: imageROM = 8'd29;
                28: imageROM = 8'd102;
                29: imageROM = 8'd63;
                30: imageROM = 8'd25;
                31: imageROM = 8'd106;
                32: imageROM = 8'd63;
                33: imageROM = 8'd21;
                34: imageROM = 8'd78;
                35: imageROM = 8'd146;
                36: imageROM = 8'd77;
                37: imageROM = 8'd63;
                38: imageROM = 8'd18;
                39: imageROM = 8'd76;
                40: imageROM = 8'd154;
                41: imageROM = 8'd74;
                42: imageROM = 8'd63;
                43: imageROM = 8'd16;
                44: imageROM = 8'd75;
                45: imageROM = 8'd158;
                46: imageROM = 8'd73;
                47: imageROM = 8'd63;
                48: imageROM = 8'd14;
                49: imageROM = 8'd73;
                50: imageROM = 8'd163;
                51: imageROM = 8'd72;
                52: imageROM = 8'd63;
                53: imageROM = 8'd12;
                54: imageROM = 8'd73;
                55: imageROM = 8'd165;
                56: imageROM = 8'd72;
                57: imageROM = 8'd63;
                58: imageROM = 8'd10;
                59: imageROM = 8'd72;
                60: imageROM = 8'd168;
                61: imageROM = 8'd72;
                62: imageROM = 8'd63;
                63: imageROM = 8'd8;
                64: imageROM = 8'd72;
                65: imageROM = 8'd171;
                66: imageROM = 8'd71;
                67: imageROM = 8'd63;
                68: imageROM = 8'd6;
                69: imageROM = 8'd71;
                70: imageROM = 8'd135;
                71: imageROM = 8'd69;
                72: imageROM = 8'd161;
                73: imageROM = 8'd71;
                74: imageROM = 8'd63;
                75: imageROM = 8'd5;
                76: imageROM = 8'd71;
                77: imageROM = 8'd135;
                78: imageROM = 8'd71;
                79: imageROM = 8'd159;
                80: imageROM = 8'd73;
                81: imageROM = 8'd63;
                82: imageROM = 8'd3;
                83: imageROM = 8'd71;
                84: imageROM = 8'd135;
                85: imageROM = 8'd73;
                86: imageROM = 8'd141;
                87: imageROM = 8'd72;
                88: imageROM = 8'd136;
                89: imageROM = 8'd74;
                90: imageROM = 8'd63;
                91: imageROM = 8'd2;
                92: imageROM = 8'd71;
                93: imageROM = 8'd136;
                94: imageROM = 8'd73;
                95: imageROM = 8'd139;
                96: imageROM = 8'd76;
                97: imageROM = 8'd134;
                98: imageROM = 8'd75;
                99: imageROM = 8'd63;
                100: imageROM = 8'd1;
                101: imageROM = 8'd70;
                102: imageROM = 8'd137;
                103: imageROM = 8'd74;
                104: imageROM = 8'd136;
                105: imageROM = 8'd79;
                106: imageROM = 8'd133;
                107: imageROM = 8'd75;
                108: imageROM = 8'd63;
                109: imageROM = 8'd70;
                110: imageROM = 8'd138;
                111: imageROM = 8'd74;
                112: imageROM = 8'd135;
                113: imageROM = 8'd81;
                114: imageROM = 8'd132;
                115: imageROM = 8'd76;
                116: imageROM = 8'd61;
                117: imageROM = 8'd71;
                118: imageROM = 8'd138;
                119: imageROM = 8'd74;
                120: imageROM = 8'd135;
                121: imageROM = 8'd82;
                122: imageROM = 8'd131;
                123: imageROM = 8'd76;
                124: imageROM = 8'd61;
                125: imageROM = 8'd70;
                126: imageROM = 8'd139;
                127: imageROM = 8'd74;
                128: imageROM = 8'd134;
                129: imageROM = 8'd84;
                130: imageROM = 8'd130;
                131: imageROM = 8'd77;
                132: imageROM = 8'd59;
                133: imageROM = 8'd70;
                134: imageROM = 8'd140;
                135: imageROM = 8'd74;
                136: imageROM = 8'd134;
                137: imageROM = 8'd70;
                138: imageROM = 8'd199;
                139: imageROM = 8'd71;
                140: imageROM = 8'd130;
                141: imageROM = 8'd77;
                142: imageROM = 8'd59;
                143: imageROM = 8'd70;
                144: imageROM = 8'd140;
                145: imageROM = 8'd74;
                146: imageROM = 8'd133;
                147: imageROM = 8'd71;
                148: imageROM = 8'd200;
                149: imageROM = 8'd71;
                150: imageROM = 8'd130;
                151: imageROM = 8'd76;
                152: imageROM = 8'd58;
                153: imageROM = 8'd70;
                154: imageROM = 8'd142;
                155: imageROM = 8'd73;
                156: imageROM = 8'd133;
                157: imageROM = 8'd70;
                158: imageROM = 8'd202;
                159: imageROM = 8'd70;
                160: imageROM = 8'd131;
                161: imageROM = 8'd69;
                162: imageROM = 8'd129;
                163: imageROM = 8'd70;
                164: imageROM = 8'd57;
                165: imageROM = 8'd70;
                166: imageROM = 8'd143;
                167: imageROM = 8'd71;
                168: imageROM = 8'd134;
                169: imageROM = 8'd70;
                170: imageROM = 8'd202;
                171: imageROM = 8'd70;
                172: imageROM = 8'd133;
                173: imageROM = 8'd66;
                174: imageROM = 8'd130;
                175: imageROM = 8'd70;
                176: imageROM = 8'd57;
                177: imageROM = 8'd70;
                178: imageROM = 8'd144;
                179: imageROM = 8'd69;
                180: imageROM = 8'd134;
                181: imageROM = 8'd70;
                182: imageROM = 8'd204;
                183: imageROM = 8'd70;
                184: imageROM = 8'd137;
                185: imageROM = 8'd70;
                186: imageROM = 8'd55;
                187: imageROM = 8'd70;
                188: imageROM = 8'd156;
                189: imageROM = 8'd70;
                190: imageROM = 8'd204;
                191: imageROM = 8'd70;
                192: imageROM = 8'd137;
                193: imageROM = 8'd70;
                194: imageROM = 8'd55;
                195: imageROM = 8'd70;
                196: imageROM = 8'd156;
                197: imageROM = 8'd70;
                198: imageROM = 8'd204;
                199: imageROM = 8'd70;
                200: imageROM = 8'd138;
                201: imageROM = 8'd70;
                202: imageROM = 8'd54;
                203: imageROM = 8'd69;
                204: imageROM = 8'd157;
                205: imageROM = 8'd70;
                206: imageROM = 8'd204;
                207: imageROM = 8'd70;
                208: imageROM = 8'd139;
                209: imageROM = 8'd69;
                210: imageROM = 8'd53;
                211: imageROM = 8'd70;
                212: imageROM = 8'd157;
                213: imageROM = 8'd70;
                214: imageROM = 8'd205;
                215: imageROM = 8'd69;
                216: imageROM = 8'd139;
                217: imageROM = 8'd70;
                218: imageROM = 8'd52;
                219: imageROM = 8'd70;
                220: imageROM = 8'd157;
                221: imageROM = 8'd70;
                222: imageROM = 8'd205;
                223: imageROM = 8'd70;
                224: imageROM = 8'd138;
                225: imageROM = 8'd70;
                226: imageROM = 8'd52;
                227: imageROM = 8'd70;
                228: imageROM = 8'd156;
                229: imageROM = 8'd71;
                230: imageROM = 8'd205;
                231: imageROM = 8'd70;
                232: imageROM = 8'd139;
                233: imageROM = 8'd69;
                234: imageROM = 8'd52;
                235: imageROM = 8'd69;
                236: imageROM = 8'd158;
                237: imageROM = 8'd70;
                238: imageROM = 8'd205;
                239: imageROM = 8'd70;
                240: imageROM = 8'd139;
                241: imageROM = 8'd70;
                242: imageROM = 8'd50;
                243: imageROM = 8'd70;
                244: imageROM = 8'd158;
                245: imageROM = 8'd70;
                246: imageROM = 8'd205;
                247: imageROM = 8'd70;
                248: imageROM = 8'd139;
                249: imageROM = 8'd70;
                250: imageROM = 8'd50;
                251: imageROM = 8'd70;
                252: imageROM = 8'd158;
                253: imageROM = 8'd70;
                254: imageROM = 8'd205;
                255: imageROM = 8'd70;
                256: imageROM = 8'd139;
                257: imageROM = 8'd70;
                258: imageROM = 8'd50;
                259: imageROM = 8'd70;
                260: imageROM = 8'd158;
                261: imageROM = 8'd70;
                262: imageROM = 8'd205;
                263: imageROM = 8'd70;
                264: imageROM = 8'd140;
                265: imageROM = 8'd69;
                266: imageROM = 8'd50;
                267: imageROM = 8'd69;
                268: imageROM = 8'd159;
                269: imageROM = 8'd70;
                270: imageROM = 8'd205;
                271: imageROM = 8'd70;
                272: imageROM = 8'd140;
                273: imageROM = 8'd70;
                274: imageROM = 8'd48;
                275: imageROM = 8'd70;
                276: imageROM = 8'd159;
                277: imageROM = 8'd70;
                278: imageROM = 8'd205;
                279: imageROM = 8'd70;
                280: imageROM = 8'd140;
                281: imageROM = 8'd70;
                282: imageROM = 8'd48;
                283: imageROM = 8'd70;
                284: imageROM = 8'd159;
                285: imageROM = 8'd70;
                286: imageROM = 8'd205;
                287: imageROM = 8'd70;
                288: imageROM = 8'd140;
                289: imageROM = 8'd70;
                290: imageROM = 8'd47;
                291: imageROM = 8'd70;
                292: imageROM = 8'd161;
                293: imageROM = 8'd70;
                294: imageROM = 8'd204;
                295: imageROM = 8'd70;
                296: imageROM = 8'd141;
                297: imageROM = 8'd69;
                298: imageROM = 8'd47;
                299: imageROM = 8'd70;
                300: imageROM = 8'd161;
                301: imageROM = 8'd70;
                302: imageROM = 8'd203;
                303: imageROM = 8'd70;
                304: imageROM = 8'd142;
                305: imageROM = 8'd69;
                306: imageROM = 8'd47;
                307: imageROM = 8'd69;
                308: imageROM = 8'd162;
                309: imageROM = 8'd70;
                310: imageROM = 8'd203;
                311: imageROM = 8'd70;
                312: imageROM = 8'd142;
                313: imageROM = 8'd69;
                314: imageROM = 8'd46;
                315: imageROM = 8'd70;
                316: imageROM = 8'd162;
                317: imageROM = 8'd70;
                318: imageROM = 8'd203;
                319: imageROM = 8'd70;
                320: imageROM = 8'd142;
                321: imageROM = 8'd69;
                322: imageROM = 8'd46;
                323: imageROM = 8'd70;
                324: imageROM = 8'd163;
                325: imageROM = 8'd69;
                326: imageROM = 8'd203;
                327: imageROM = 8'd70;
                328: imageROM = 8'd142;
                329: imageROM = 8'd69;
                330: imageROM = 8'd45;
                331: imageROM = 8'd70;
                332: imageROM = 8'd164;
                333: imageROM = 8'd70;
                334: imageROM = 8'd201;
                335: imageROM = 8'd70;
                336: imageROM = 8'd143;
                337: imageROM = 8'd69;
                338: imageROM = 8'd45;
                339: imageROM = 8'd70;
                340: imageROM = 8'd164;
                341: imageROM = 8'd70;
                342: imageROM = 8'd201;
                343: imageROM = 8'd70;
                344: imageROM = 8'd142;
                345: imageROM = 8'd70;
                346: imageROM = 8'd44;
                347: imageROM = 8'd71;
                348: imageROM = 8'd165;
                349: imageROM = 8'd70;
                350: imageROM = 8'd199;
                351: imageROM = 8'd71;
                352: imageROM = 8'd142;
                353: imageROM = 8'd70;
                354: imageROM = 8'd44;
                355: imageROM = 8'd70;
                356: imageROM = 8'd166;
                357: imageROM = 8'd70;
                358: imageROM = 8'd198;
                359: imageROM = 8'd71;
                360: imageROM = 8'd143;
                361: imageROM = 8'd70;
                362: imageROM = 8'd43;
                363: imageROM = 8'd71;
                364: imageROM = 8'd166;
                365: imageROM = 8'd71;
                366: imageROM = 8'd197;
                367: imageROM = 8'd71;
                368: imageROM = 8'd143;
                369: imageROM = 8'd70;
                370: imageROM = 8'd43;
                371: imageROM = 8'd71;
                372: imageROM = 8'd167;
                373: imageROM = 8'd71;
                374: imageROM = 8'd195;
                375: imageROM = 8'd71;
                376: imageROM = 8'd144;
                377: imageROM = 8'd69;
                378: imageROM = 8'd43;
                379: imageROM = 8'd72;
                380: imageROM = 8'd168;
                381: imageROM = 8'd70;
                382: imageROM = 8'd195;
                383: imageROM = 8'd70;
                384: imageROM = 8'd144;
                385: imageROM = 8'd70;
                386: imageROM = 8'd43;
                387: imageROM = 8'd72;
                388: imageROM = 8'd168;
                389: imageROM = 8'd71;
                390: imageROM = 8'd193;
                391: imageROM = 8'd71;
                392: imageROM = 8'd144;
                393: imageROM = 8'd70;
                394: imageROM = 8'd42;
                395: imageROM = 8'd73;
                396: imageROM = 8'd169;
                397: imageROM = 8'd77;
                398: imageROM = 8'd145;
                399: imageROM = 8'd70;
                400: imageROM = 8'd41;
                401: imageROM = 8'd74;
                402: imageROM = 8'd170;
                403: imageROM = 8'd76;
                404: imageROM = 8'd145;
                405: imageROM = 8'd69;
                406: imageROM = 8'd42;
                407: imageROM = 8'd75;
                408: imageROM = 8'd170;
                409: imageROM = 8'd74;
                410: imageROM = 8'd145;
                411: imageROM = 8'd70;
                412: imageROM = 8'd41;
                413: imageROM = 8'd76;
                414: imageROM = 8'd170;
                415: imageROM = 8'd73;
                416: imageROM = 8'd146;
                417: imageROM = 8'd70;
                418: imageROM = 8'd41;
                419: imageROM = 8'd76;
                420: imageROM = 8'd171;
                421: imageROM = 8'd72;
                422: imageROM = 8'd146;
                423: imageROM = 8'd69;
                424: imageROM = 8'd41;
                425: imageROM = 8'd70;
                426: imageROM = 8'd130;
                427: imageROM = 8'd70;
                428: imageROM = 8'd171;
                429: imageROM = 8'd70;
                430: imageROM = 8'd146;
                431: imageROM = 8'd70;
                432: imageROM = 8'd40;
                433: imageROM = 8'd71;
                434: imageROM = 8'd130;
                435: imageROM = 8'd70;
                436: imageROM = 8'd171;
                437: imageROM = 8'd70;
                438: imageROM = 8'd146;
                439: imageROM = 8'd70;
                440: imageROM = 8'd39;
                441: imageROM = 8'd71;
                442: imageROM = 8'd132;
                443: imageROM = 8'd70;
                444: imageROM = 8'd171;
                445: imageROM = 8'd68;
                446: imageROM = 8'd146;
                447: imageROM = 8'd70;
                448: imageROM = 8'd40;
                449: imageROM = 8'd70;
                450: imageROM = 8'd133;
                451: imageROM = 8'd70;
                452: imageROM = 8'd172;
                453: imageROM = 8'd67;
                454: imageROM = 8'd146;
                455: imageROM = 8'd70;
                456: imageROM = 8'd39;
                457: imageROM = 8'd71;
                458: imageROM = 8'd134;
                459: imageROM = 8'd70;
                460: imageROM = 8'd191;
                461: imageROM = 8'd129;
                462: imageROM = 8'd70;
                463: imageROM = 8'd38;
                464: imageROM = 8'd71;
                465: imageROM = 8'd135;
                466: imageROM = 8'd71;
                467: imageROM = 8'd190;
                468: imageROM = 8'd70;
                469: imageROM = 8'd38;
                470: imageROM = 8'd71;
                471: imageROM = 8'd137;
                472: imageROM = 8'd70;
                473: imageROM = 8'd190;
                474: imageROM = 8'd70;
                475: imageROM = 8'd37;
                476: imageROM = 8'd71;
                477: imageROM = 8'd139;
                478: imageROM = 8'd70;
                479: imageROM = 8'd189;
                480: imageROM = 8'd69;
                481: imageROM = 8'd37;
                482: imageROM = 8'd71;
                483: imageROM = 8'd140;
                484: imageROM = 8'd71;
                485: imageROM = 8'd187;
                486: imageROM = 8'd70;
                487: imageROM = 8'd36;
                488: imageROM = 8'd72;
                489: imageROM = 8'd141;
                490: imageROM = 8'd71;
                491: imageROM = 8'd186;
                492: imageROM = 8'd70;
                493: imageROM = 8'd35;
                494: imageROM = 8'd72;
                495: imageROM = 8'd143;
                496: imageROM = 8'd71;
                497: imageROM = 8'd185;
                498: imageROM = 8'd69;
                499: imageROM = 8'd35;
                500: imageROM = 8'd72;
                501: imageROM = 8'd145;
                502: imageROM = 8'd72;
                503: imageROM = 8'd182;
                504: imageROM = 8'd70;
                505: imageROM = 8'd35;
                506: imageROM = 8'd71;
                507: imageROM = 8'd147;
                508: imageROM = 8'd72;
                509: imageROM = 8'd181;
                510: imageROM = 8'd70;
                511: imageROM = 8'd34;
                512: imageROM = 8'd71;
                513: imageROM = 8'd149;
                514: imageROM = 8'd73;
                515: imageROM = 8'd179;
                516: imageROM = 8'd69;
                517: imageROM = 8'd34;
                518: imageROM = 8'd71;
                519: imageROM = 8'd151;
                520: imageROM = 8'd74;
                521: imageROM = 8'd176;
                522: imageROM = 8'd70;
                523: imageROM = 8'd33;
                524: imageROM = 8'd71;
                525: imageROM = 8'd153;
                526: imageROM = 8'd77;
                527: imageROM = 8'd172;
                528: imageROM = 8'd70;
                529: imageROM = 8'd32;
                530: imageROM = 8'd71;
                531: imageROM = 8'd156;
                532: imageROM = 8'd82;
                533: imageROM = 8'd165;
                534: imageROM = 8'd70;
                535: imageROM = 8'd32;
                536: imageROM = 8'd71;
                537: imageROM = 8'd157;
                538: imageROM = 8'd81;
                539: imageROM = 8'd165;
                540: imageROM = 8'd70;
                541: imageROM = 8'd31;
                542: imageROM = 8'd71;
                543: imageROM = 8'd160;
                544: imageROM = 8'd79;
                545: imageROM = 8'd165;
                546: imageROM = 8'd70;
                547: imageROM = 8'd30;
                548: imageROM = 8'd71;
                549: imageROM = 8'd164;
                550: imageROM = 8'd76;
                551: imageROM = 8'd165;
                552: imageROM = 8'd70;
                553: imageROM = 8'd29;
                554: imageROM = 8'd71;
                555: imageROM = 8'd167;
                556: imageROM = 8'd74;
                557: imageROM = 8'd165;
                558: imageROM = 8'd69;
                559: imageROM = 8'd29;
                560: imageROM = 8'd71;
                561: imageROM = 8'd174;
                562: imageROM = 8'd66;
                563: imageROM = 8'd167;
                564: imageROM = 8'd69;
                565: imageROM = 8'd28;
                566: imageROM = 8'd71;
                567: imageROM = 8'd191;
                568: imageROM = 8'd153;
                569: imageROM = 8'd70;
                570: imageROM = 8'd26;
                571: imageROM = 8'd71;
                572: imageROM = 8'd191;
                573: imageROM = 8'd154;
                574: imageROM = 8'd70;
                575: imageROM = 8'd25;
                576: imageROM = 8'd71;
                577: imageROM = 8'd191;
                578: imageROM = 8'd155;
                579: imageROM = 8'd70;
                580: imageROM = 8'd24;
                581: imageROM = 8'd71;
                582: imageROM = 8'd191;
                583: imageROM = 8'd156;
                584: imageROM = 8'd70;
                585: imageROM = 8'd23;
                586: imageROM = 8'd71;
                587: imageROM = 8'd191;
                588: imageROM = 8'd157;
                589: imageROM = 8'd70;
                590: imageROM = 8'd22;
                591: imageROM = 8'd71;
                592: imageROM = 8'd191;
                593: imageROM = 8'd158;
                594: imageROM = 8'd70;
                595: imageROM = 8'd21;
                596: imageROM = 8'd71;
                597: imageROM = 8'd191;
                598: imageROM = 8'd160;
                599: imageROM = 8'd69;
                600: imageROM = 8'd20;
                601: imageROM = 8'd71;
                602: imageROM = 8'd191;
                603: imageROM = 8'd161;
                604: imageROM = 8'd70;
                605: imageROM = 8'd18;
                606: imageROM = 8'd71;
                607: imageROM = 8'd191;
                608: imageROM = 8'd162;
                609: imageROM = 8'd70;
                610: imageROM = 8'd18;
                611: imageROM = 8'd70;
                612: imageROM = 8'd191;
                613: imageROM = 8'd163;
                614: imageROM = 8'd70;
                615: imageROM = 8'd17;
                616: imageROM = 8'd70;
                617: imageROM = 8'd191;
                618: imageROM = 8'd165;
                619: imageROM = 8'd69;
                620: imageROM = 8'd17;
                621: imageROM = 8'd70;
                622: imageROM = 8'd191;
                623: imageROM = 8'd165;
                624: imageROM = 8'd70;
                625: imageROM = 8'd16;
                626: imageROM = 8'd69;
                627: imageROM = 8'd191;
                628: imageROM = 8'd167;
                629: imageROM = 8'd69;
            // r02.bmp
                630: imageROM = 8'd57;
                631: imageROM = 8'd76;
                632: imageROM = 8'd63;
                633: imageROM = 8'd50;
                634: imageROM = 8'd83;
                635: imageROM = 8'd63;
                636: imageROM = 8'd43;
                637: imageROM = 8'd89;
                638: imageROM = 8'd63;
                639: imageROM = 8'd38;
                640: imageROM = 8'd92;
                641: imageROM = 8'd63;
                642: imageROM = 8'd35;
                643: imageROM = 8'd96;
                644: imageROM = 8'd63;
                645: imageROM = 8'd32;
                646: imageROM = 8'd98;
                647: imageROM = 8'd63;
                648: imageROM = 8'd29;
                649: imageROM = 8'd77;
                650: imageROM = 8'd141;
                651: imageROM = 8'd75;
                652: imageROM = 8'd63;
                653: imageROM = 8'd27;
                654: imageROM = 8'd75;
                655: imageROM = 8'd147;
                656: imageROM = 8'd73;
                657: imageROM = 8'd63;
                658: imageROM = 8'd24;
                659: imageROM = 8'd75;
                660: imageROM = 8'd151;
                661: imageROM = 8'd72;
                662: imageROM = 8'd63;
                663: imageROM = 8'd22;
                664: imageROM = 8'd74;
                665: imageROM = 8'd154;
                666: imageROM = 8'd72;
                667: imageROM = 8'd63;
                668: imageROM = 8'd20;
                669: imageROM = 8'd73;
                670: imageROM = 8'd158;
                671: imageROM = 8'd71;
                672: imageROM = 8'd63;
                673: imageROM = 8'd18;
                674: imageROM = 8'd73;
                675: imageROM = 8'd160;
                676: imageROM = 8'd71;
                677: imageROM = 8'd63;
                678: imageROM = 8'd16;
                679: imageROM = 8'd72;
                680: imageROM = 8'd163;
                681: imageROM = 8'd71;
                682: imageROM = 8'd63;
                683: imageROM = 8'd14;
                684: imageROM = 8'd75;
                685: imageROM = 8'd162;
                686: imageROM = 8'd71;
                687: imageROM = 8'd63;
                688: imageROM = 8'd12;
                689: imageROM = 8'd78;
                690: imageROM = 8'd160;
                691: imageROM = 8'd71;
                692: imageROM = 8'd63;
                693: imageROM = 8'd11;
                694: imageROM = 8'd79;
                695: imageROM = 8'd158;
                696: imageROM = 8'd74;
                697: imageROM = 8'd63;
                698: imageROM = 8'd9;
                699: imageROM = 8'd81;
                700: imageROM = 8'd157;
                701: imageROM = 8'd75;
                702: imageROM = 8'd63;
                703: imageROM = 8'd8;
                704: imageROM = 8'd81;
                705: imageROM = 8'd144;
                706: imageROM = 8'd68;
                707: imageROM = 8'd136;
                708: imageROM = 8'd77;
                709: imageROM = 8'd63;
                710: imageROM = 8'd6;
                711: imageROM = 8'd71;
                712: imageROM = 8'd130;
                713: imageROM = 8'd74;
                714: imageROM = 8'd139;
                715: imageROM = 8'd75;
                716: imageROM = 8'd133;
                717: imageROM = 8'd77;
                718: imageROM = 8'd63;
                719: imageROM = 8'd5;
                720: imageROM = 8'd71;
                721: imageROM = 8'd131;
                722: imageROM = 8'd74;
                723: imageROM = 8'd138;
                724: imageROM = 8'd77;
                725: imageROM = 8'd132;
                726: imageROM = 8'd78;
                727: imageROM = 8'd63;
                728: imageROM = 8'd4;
                729: imageROM = 8'd71;
                730: imageROM = 8'd131;
                731: imageROM = 8'd74;
                732: imageROM = 8'd137;
                733: imageROM = 8'd79;
                734: imageROM = 8'd131;
                735: imageROM = 8'd79;
                736: imageROM = 8'd63;
                737: imageROM = 8'd2;
                738: imageROM = 8'd71;
                739: imageROM = 8'd132;
                740: imageROM = 8'd74;
                741: imageROM = 8'd136;
                742: imageROM = 8'd81;
                743: imageROM = 8'd130;
                744: imageROM = 8'd79;
                745: imageROM = 8'd63;
                746: imageROM = 8'd2;
                747: imageROM = 8'd70;
                748: imageROM = 8'd133;
                749: imageROM = 8'd74;
                750: imageROM = 8'd135;
                751: imageROM = 8'd83;
                752: imageROM = 8'd130;
                753: imageROM = 8'd71;
                754: imageROM = 8'd129;
                755: imageROM = 8'd71;
                756: imageROM = 8'd63;
                757: imageROM = 8'd71;
                758: imageROM = 8'd133;
                759: imageROM = 8'd74;
                760: imageROM = 8'd135;
                761: imageROM = 8'd71;
                762: imageROM = 8'd197;
                763: imageROM = 8'd72;
                764: imageROM = 8'd129;
                765: imageROM = 8'd71;
                766: imageROM = 8'd130;
                767: imageROM = 8'd70;
                768: imageROM = 8'd63;
                769: imageROM = 8'd70;
                770: imageROM = 8'd135;
                771: imageROM = 8'd72;
                772: imageROM = 8'd135;
                773: imageROM = 8'd71;
                774: imageROM = 8'd200;
                775: imageROM = 8'd70;
                776: imageROM = 8'd131;
                777: imageROM = 8'd68;
                778: imageROM = 8'd132;
                779: imageROM = 8'd70;
                780: imageROM = 8'd61;
                781: imageROM = 8'd70;
                782: imageROM = 8'd137;
                783: imageROM = 8'd71;
                784: imageROM = 8'd135;
                785: imageROM = 8'd70;
                786: imageROM = 8'd201;
                787: imageROM = 8'd71;
                788: imageROM = 8'd138;
                789: imageROM = 8'd71;
                790: imageROM = 8'd60;
                791: imageROM = 8'd70;
                792: imageROM = 8'd138;
                793: imageROM = 8'd68;
                794: imageROM = 8'd137;
                795: imageROM = 8'd69;
                796: imageROM = 8'd203;
                797: imageROM = 8'd70;
                798: imageROM = 8'd139;
                799: imageROM = 8'd70;
                800: imageROM = 8'd59;
                801: imageROM = 8'd71;
                802: imageROM = 8'd150;
                803: imageROM = 8'd70;
                804: imageROM = 8'd203;
                805: imageROM = 8'd70;
                806: imageROM = 8'd139;
                807: imageROM = 8'd71;
                808: imageROM = 8'd58;
                809: imageROM = 8'd70;
                810: imageROM = 8'd151;
                811: imageROM = 8'd70;
                812: imageROM = 8'd204;
                813: imageROM = 8'd70;
                814: imageROM = 8'd139;
                815: imageROM = 8'd70;
                816: imageROM = 8'd58;
                817: imageROM = 8'd70;
                818: imageROM = 8'd151;
                819: imageROM = 8'd70;
                820: imageROM = 8'd204;
                821: imageROM = 8'd70;
                822: imageROM = 8'd139;
                823: imageROM = 8'd71;
                824: imageROM = 8'd56;
                825: imageROM = 8'd70;
                826: imageROM = 8'd152;
                827: imageROM = 8'd69;
                828: imageROM = 8'd205;
                829: imageROM = 8'd70;
                830: imageROM = 8'd140;
                831: imageROM = 8'd70;
                832: imageROM = 8'd56;
                833: imageROM = 8'd70;
                834: imageROM = 8'd152;
                835: imageROM = 8'd69;
                836: imageROM = 8'd205;
                837: imageROM = 8'd70;
                838: imageROM = 8'd140;
                839: imageROM = 8'd70;
                840: imageROM = 8'd56;
                841: imageROM = 8'd70;
                842: imageROM = 8'd152;
                843: imageROM = 8'd69;
                844: imageROM = 8'd206;
                845: imageROM = 8'd69;
                846: imageROM = 8'd140;
                847: imageROM = 8'd70;
                848: imageROM = 8'd56;
                849: imageROM = 8'd69;
                850: imageROM = 8'd152;
                851: imageROM = 8'd70;
                852: imageROM = 8'd206;
                853: imageROM = 8'd69;
                854: imageROM = 8'd141;
                855: imageROM = 8'd70;
                856: imageROM = 8'd54;
                857: imageROM = 8'd70;
                858: imageROM = 8'd152;
                859: imageROM = 8'd70;
                860: imageROM = 8'd206;
                861: imageROM = 8'd69;
                862: imageROM = 8'd141;
                863: imageROM = 8'd70;
                864: imageROM = 8'd54;
                865: imageROM = 8'd70;
                866: imageROM = 8'd152;
                867: imageROM = 8'd70;
                868: imageROM = 8'd206;
                869: imageROM = 8'd70;
                870: imageROM = 8'd140;
                871: imageROM = 8'd70;
                872: imageROM = 8'd54;
                873: imageROM = 8'd70;
                874: imageROM = 8'd153;
                875: imageROM = 8'd69;
                876: imageROM = 8'd206;
                877: imageROM = 8'd70;
                878: imageROM = 8'd140;
                879: imageROM = 8'd70;
                880: imageROM = 8'd54;
                881: imageROM = 8'd70;
                882: imageROM = 8'd153;
                883: imageROM = 8'd69;
                884: imageROM = 8'd206;
                885: imageROM = 8'd70;
                886: imageROM = 8'd140;
                887: imageROM = 8'd70;
                888: imageROM = 8'd54;
                889: imageROM = 8'd69;
                890: imageROM = 8'd154;
                891: imageROM = 8'd69;
                892: imageROM = 8'd206;
                893: imageROM = 8'd70;
                894: imageROM = 8'd140;
                895: imageROM = 8'd70;
                896: imageROM = 8'd53;
                897: imageROM = 8'd70;
                898: imageROM = 8'd154;
                899: imageROM = 8'd70;
                900: imageROM = 8'd205;
                901: imageROM = 8'd70;
                902: imageROM = 8'd141;
                903: imageROM = 8'd69;
                904: imageROM = 8'd53;
                905: imageROM = 8'd70;
                906: imageROM = 8'd154;
                907: imageROM = 8'd70;
                908: imageROM = 8'd205;
                909: imageROM = 8'd69;
                910: imageROM = 8'd142;
                911: imageROM = 8'd70;
                912: imageROM = 8'd52;
                913: imageROM = 8'd70;
                914: imageROM = 8'd154;
                915: imageROM = 8'd70;
                916: imageROM = 8'd205;
                917: imageROM = 8'd69;
                918: imageROM = 8'd142;
                919: imageROM = 8'd70;
                920: imageROM = 8'd52;
                921: imageROM = 8'd70;
                922: imageROM = 8'd154;
                923: imageROM = 8'd70;
                924: imageROM = 8'd204;
                925: imageROM = 8'd70;
                926: imageROM = 8'd142;
                927: imageROM = 8'd70;
                928: imageROM = 8'd52;
                929: imageROM = 8'd69;
                930: imageROM = 8'd156;
                931: imageROM = 8'd69;
                932: imageROM = 8'd204;
                933: imageROM = 8'd70;
                934: imageROM = 8'd142;
                935: imageROM = 8'd70;
                936: imageROM = 8'd51;
                937: imageROM = 8'd70;
                938: imageROM = 8'd156;
                939: imageROM = 8'd70;
                940: imageROM = 8'd203;
                941: imageROM = 8'd70;
                942: imageROM = 8'd142;
                943: imageROM = 8'd70;
                944: imageROM = 8'd51;
                945: imageROM = 8'd70;
                946: imageROM = 8'd156;
                947: imageROM = 8'd70;
                948: imageROM = 8'd203;
                949: imageROM = 8'd70;
                950: imageROM = 8'd142;
                951: imageROM = 8'd70;
                952: imageROM = 8'd51;
                953: imageROM = 8'd70;
                954: imageROM = 8'd156;
                955: imageROM = 8'd70;
                956: imageROM = 8'd202;
                957: imageROM = 8'd70;
                958: imageROM = 8'd143;
                959: imageROM = 8'd70;
                960: imageROM = 8'd51;
                961: imageROM = 8'd70;
                962: imageROM = 8'd157;
                963: imageROM = 8'd70;
                964: imageROM = 8'd201;
                965: imageROM = 8'd70;
                966: imageROM = 8'd143;
                967: imageROM = 8'd70;
                968: imageROM = 8'd51;
                969: imageROM = 8'd70;
                970: imageROM = 8'd157;
                971: imageROM = 8'd70;
                972: imageROM = 8'd200;
                973: imageROM = 8'd71;
                974: imageROM = 8'd143;
                975: imageROM = 8'd70;
                976: imageROM = 8'd50;
                977: imageROM = 8'd71;
                978: imageROM = 8'd157;
                979: imageROM = 8'd71;
                980: imageROM = 8'd199;
                981: imageROM = 8'd70;
                982: imageROM = 8'd144;
                983: imageROM = 8'd70;
                984: imageROM = 8'd50;
                985: imageROM = 8'd70;
                986: imageROM = 8'd159;
                987: imageROM = 8'd70;
                988: imageROM = 8'd198;
                989: imageROM = 8'd71;
                990: imageROM = 8'd144;
                991: imageROM = 8'd70;
                992: imageROM = 8'd50;
                993: imageROM = 8'd70;
                994: imageROM = 8'd159;
                995: imageROM = 8'd71;
                996: imageROM = 8'd196;
                997: imageROM = 8'd71;
                998: imageROM = 8'd145;
                999: imageROM = 8'd70;
                1000: imageROM = 8'd50;
                1001: imageROM = 8'd70;
                1002: imageROM = 8'd160;
                1003: imageROM = 8'd71;
                1004: imageROM = 8'd195;
                1005: imageROM = 8'd70;
                1006: imageROM = 8'd146;
                1007: imageROM = 8'd70;
                1008: imageROM = 8'd50;
                1009: imageROM = 8'd70;
                1010: imageROM = 8'd161;
                1011: imageROM = 8'd71;
                1012: imageROM = 8'd193;
                1013: imageROM = 8'd71;
                1014: imageROM = 8'd147;
                1015: imageROM = 8'd69;
                1016: imageROM = 8'd50;
                1017: imageROM = 8'd70;
                1018: imageROM = 8'd161;
                1019: imageROM = 8'd71;
                1020: imageROM = 8'd193;
                1021: imageROM = 8'd70;
                1022: imageROM = 8'd148;
                1023: imageROM = 8'd69;
                1024: imageROM = 8'd50;
                1025: imageROM = 8'd70;
                1026: imageROM = 8'd162;
                1027: imageROM = 8'd77;
                1028: imageROM = 8'd148;
                1029: imageROM = 8'd69;
                1030: imageROM = 8'd50;
                1031: imageROM = 8'd70;
                1032: imageROM = 8'd163;
                1033: imageROM = 8'd75;
                1034: imageROM = 8'd149;
                1035: imageROM = 8'd69;
                1036: imageROM = 8'd50;
                1037: imageROM = 8'd71;
                1038: imageROM = 8'd162;
                1039: imageROM = 8'd74;
                1040: imageROM = 8'd150;
                1041: imageROM = 8'd70;
                1042: imageROM = 8'd48;
                1043: imageROM = 8'd72;
                1044: imageROM = 8'd163;
                1045: imageROM = 8'd73;
                1046: imageROM = 8'd150;
                1047: imageROM = 8'd69;
                1048: imageROM = 8'd49;
                1049: imageROM = 8'd72;
                1050: imageROM = 8'd164;
                1051: imageROM = 8'd71;
                1052: imageROM = 8'd151;
                1053: imageROM = 8'd69;
                1054: imageROM = 8'd49;
                1055: imageROM = 8'd73;
                1056: imageROM = 8'd164;
                1057: imageROM = 8'd70;
                1058: imageROM = 8'd151;
                1059: imageROM = 8'd70;
                1060: imageROM = 8'd48;
                1061: imageROM = 8'd73;
                1062: imageROM = 8'd165;
                1063: imageROM = 8'd68;
                1064: imageROM = 8'd152;
                1065: imageROM = 8'd70;
                1066: imageROM = 8'd48;
                1067: imageROM = 8'd73;
                1068: imageROM = 8'd165;
                1069: imageROM = 8'd68;
                1070: imageROM = 8'd152;
                1071: imageROM = 8'd70;
                1072: imageROM = 8'd48;
                1073: imageROM = 8'd74;
                1074: imageROM = 8'd165;
                1075: imageROM = 8'd66;
                1076: imageROM = 8'd153;
                1077: imageROM = 8'd70;
                1078: imageROM = 8'd48;
                1079: imageROM = 8'd75;
                1080: imageROM = 8'd191;
                1081: imageROM = 8'd70;
                1082: imageROM = 8'd47;
                1083: imageROM = 8'd76;
                1084: imageROM = 8'd191;
                1085: imageROM = 8'd129;
                1086: imageROM = 8'd69;
                1087: imageROM = 8'd47;
                1088: imageROM = 8'd77;
                1089: imageROM = 8'd191;
                1090: imageROM = 8'd70;
                1091: imageROM = 8'd46;
                1092: imageROM = 8'd70;
                1093: imageROM = 8'd129;
                1094: imageROM = 8'd71;
                1095: imageROM = 8'd190;
                1096: imageROM = 8'd70;
                1097: imageROM = 8'd46;
                1098: imageROM = 8'd70;
                1099: imageROM = 8'd130;
                1100: imageROM = 8'd71;
                1101: imageROM = 8'd190;
                1102: imageROM = 8'd70;
                1103: imageROM = 8'd45;
                1104: imageROM = 8'd69;
                1105: imageROM = 8'd132;
                1106: imageROM = 8'd71;
                1107: imageROM = 8'd189;
                1108: imageROM = 8'd70;
                1109: imageROM = 8'd44;
                1110: imageROM = 8'd70;
                1111: imageROM = 8'd132;
                1112: imageROM = 8'd72;
                1113: imageROM = 8'd188;
                1114: imageROM = 8'd71;
                1115: imageROM = 8'd43;
                1116: imageROM = 8'd70;
                1117: imageROM = 8'd133;
                1118: imageROM = 8'd73;
                1119: imageROM = 8'd187;
                1120: imageROM = 8'd70;
                1121: imageROM = 8'd43;
                1122: imageROM = 8'd70;
                1123: imageROM = 8'd135;
                1124: imageROM = 8'd72;
                1125: imageROM = 8'd186;
                1126: imageROM = 8'd71;
                1127: imageROM = 8'd41;
                1128: imageROM = 8'd70;
                1129: imageROM = 8'd137;
                1130: imageROM = 8'd73;
                1131: imageROM = 8'd185;
                1132: imageROM = 8'd70;
                1133: imageROM = 8'd41;
                1134: imageROM = 8'd70;
                1135: imageROM = 8'd138;
                1136: imageROM = 8'd74;
                1137: imageROM = 8'd183;
                1138: imageROM = 8'd71;
                1139: imageROM = 8'd39;
                1140: imageROM = 8'd71;
                1141: imageROM = 8'd139;
                1142: imageROM = 8'd77;
                1143: imageROM = 8'd180;
                1144: imageROM = 8'd70;
                1145: imageROM = 8'd38;
                1146: imageROM = 8'd71;
                1147: imageROM = 8'd141;
                1148: imageROM = 8'd83;
                1149: imageROM = 8'd173;
                1150: imageROM = 8'd71;
                1151: imageROM = 8'd36;
                1152: imageROM = 8'd71;
                1153: imageROM = 8'd144;
                1154: imageROM = 8'd81;
                1155: imageROM = 8'd174;
                1156: imageROM = 8'd70;
                1157: imageROM = 8'd35;
                1158: imageROM = 8'd72;
                1159: imageROM = 8'd146;
                1160: imageROM = 8'd79;
                1161: imageROM = 8'd174;
                1162: imageROM = 8'd71;
                1163: imageROM = 8'd33;
                1164: imageROM = 8'd72;
                1165: imageROM = 8'd149;
                1166: imageROM = 8'd77;
                1167: imageROM = 8'd175;
                1168: imageROM = 8'd71;
                1169: imageROM = 8'd31;
                1170: imageROM = 8'd72;
                1171: imageROM = 8'd152;
                1172: imageROM = 8'd75;
                1173: imageROM = 8'd176;
                1174: imageROM = 8'd70;
                1175: imageROM = 8'd30;
                1176: imageROM = 8'd72;
                1177: imageROM = 8'd159;
                1178: imageROM = 8'd67;
                1179: imageROM = 8'd178;
                1180: imageROM = 8'd71;
                1181: imageROM = 8'd28;
                1182: imageROM = 8'd72;
                1183: imageROM = 8'd191;
                1184: imageROM = 8'd151;
                1185: imageROM = 8'd71;
                1186: imageROM = 8'd26;
                1187: imageROM = 8'd72;
                1188: imageROM = 8'd191;
                1189: imageROM = 8'd152;
                1190: imageROM = 8'd71;
                1191: imageROM = 8'd25;
                1192: imageROM = 8'd72;
                1193: imageROM = 8'd191;
                1194: imageROM = 8'd154;
                1195: imageROM = 8'd71;
                1196: imageROM = 8'd23;
                1197: imageROM = 8'd72;
                1198: imageROM = 8'd191;
                1199: imageROM = 8'd156;
                1200: imageROM = 8'd70;
                1201: imageROM = 8'd22;
                1202: imageROM = 8'd72;
                1203: imageROM = 8'd191;
                1204: imageROM = 8'd157;
                1205: imageROM = 8'd71;
                1206: imageROM = 8'd20;
                1207: imageROM = 8'd72;
                1208: imageROM = 8'd191;
                1209: imageROM = 8'd159;
                1210: imageROM = 8'd70;
                1211: imageROM = 8'd19;
                1212: imageROM = 8'd72;
                1213: imageROM = 8'd191;
                1214: imageROM = 8'd160;
                1215: imageROM = 8'd70;
                1216: imageROM = 8'd18;
                1217: imageROM = 8'd72;
                1218: imageROM = 8'd191;
                1219: imageROM = 8'd162;
                1220: imageROM = 8'd70;
                1221: imageROM = 8'd17;
                1222: imageROM = 8'd71;
                1223: imageROM = 8'd191;
                1224: imageROM = 8'd163;
                1225: imageROM = 8'd70;
                1226: imageROM = 8'd16;
                1227: imageROM = 8'd71;
                1228: imageROM = 8'd191;
                1229: imageROM = 8'd164;
                1230: imageROM = 8'd70;
                1231: imageROM = 8'd16;
                1232: imageROM = 8'd70;
                1233: imageROM = 8'd191;
                1234: imageROM = 8'd166;
                1235: imageROM = 8'd70;
                1236: imageROM = 8'd14;
                1237: imageROM = 8'd71;
                1238: imageROM = 8'd191;
                1239: imageROM = 8'd166;
                1240: imageROM = 8'd70;
                1241: imageROM = 8'd14;
                1242: imageROM = 8'd70;
                1243: imageROM = 8'd191;
                1244: imageROM = 8'd167;
                1245: imageROM = 8'd70;
                1246: imageROM = 8'd14;
                1247: imageROM = 8'd70;
                1248: imageROM = 8'd191;
                1249: imageROM = 8'd167;
                1250: imageROM = 8'd70;
                1251: imageROM = 8'd14;
                1252: imageROM = 8'd70;
                1253: imageROM = 8'd191;
                1254: imageROM = 8'd168;
                1255: imageROM = 8'd70;
                1256: imageROM = 8'd12;
                1257: imageROM = 8'd70;
                1258: imageROM = 8'd191;
                1259: imageROM = 8'd169;
                1260: imageROM = 8'd70;
                1261: imageROM = 8'd12;
                1262: imageROM = 8'd70;
                1263: imageROM = 8'd191;
                1264: imageROM = 8'd169;
                1265: imageROM = 8'd69;
            // r03.bmp
                1266: imageROM = 8'd63;
                1267: imageROM = 8'd63;
                1268: imageROM = 8'd63;
                1269: imageROM = 8'd63;
                1270: imageROM = 8'd63;
                1271: imageROM = 8'd63;
                1272: imageROM = 8'd43;
                1273: imageROM = 8'd81;
                1274: imageROM = 8'd63;
                1275: imageROM = 8'd44;
                1276: imageROM = 8'd89;
                1277: imageROM = 8'd63;
                1278: imageROM = 8'd37;
                1279: imageROM = 8'd95;
                1280: imageROM = 8'd63;
                1281: imageROM = 8'd32;
                1282: imageROM = 8'd99;
                1283: imageROM = 8'd63;
                1284: imageROM = 8'd28;
                1285: imageROM = 8'd102;
                1286: imageROM = 8'd63;
                1287: imageROM = 8'd25;
                1288: imageROM = 8'd105;
                1289: imageROM = 8'd63;
                1290: imageROM = 8'd23;
                1291: imageROM = 8'd76;
                1292: imageROM = 8'd149;
                1293: imageROM = 8'd75;
                1294: imageROM = 8'd63;
                1295: imageROM = 8'd20;
                1296: imageROM = 8'd74;
                1297: imageROM = 8'd155;
                1298: imageROM = 8'd72;
                1299: imageROM = 8'd63;
                1300: imageROM = 8'd19;
                1301: imageROM = 8'd73;
                1302: imageROM = 8'd158;
                1303: imageROM = 8'd72;
                1304: imageROM = 8'd63;
                1305: imageROM = 8'd17;
                1306: imageROM = 8'd72;
                1307: imageROM = 8'd162;
                1308: imageROM = 8'd71;
                1309: imageROM = 8'd63;
                1310: imageROM = 8'd15;
                1311: imageROM = 8'd72;
                1312: imageROM = 8'd164;
                1313: imageROM = 8'd71;
                1314: imageROM = 8'd63;
                1315: imageROM = 8'd13;
                1316: imageROM = 8'd71;
                1317: imageROM = 8'd167;
                1318: imageROM = 8'd71;
                1319: imageROM = 8'd63;
                1320: imageROM = 8'd11;
                1321: imageROM = 8'd71;
                1322: imageROM = 8'd155;
                1323: imageROM = 8'd68;
                1324: imageROM = 8'd137;
                1325: imageROM = 8'd71;
                1326: imageROM = 8'd63;
                1327: imageROM = 8'd10;
                1328: imageROM = 8'd71;
                1329: imageROM = 8'd134;
                1330: imageROM = 8'd69;
                1331: imageROM = 8'd142;
                1332: imageROM = 8'd74;
                1333: imageROM = 8'd135;
                1334: imageROM = 8'd71;
                1335: imageROM = 8'd63;
                1336: imageROM = 8'd8;
                1337: imageROM = 8'd71;
                1338: imageROM = 8'd133;
                1339: imageROM = 8'd72;
                1340: imageROM = 8'd140;
                1341: imageROM = 8'd76;
                1342: imageROM = 8'd135;
                1343: imageROM = 8'd70;
                1344: imageROM = 8'd63;
                1345: imageROM = 8'd8;
                1346: imageROM = 8'd70;
                1347: imageROM = 8'd134;
                1348: imageROM = 8'd72;
                1349: imageROM = 8'd139;
                1350: imageROM = 8'd79;
                1351: imageROM = 8'd132;
                1352: imageROM = 8'd72;
                1353: imageROM = 8'd63;
                1354: imageROM = 8'd6;
                1355: imageROM = 8'd71;
                1356: imageROM = 8'd133;
                1357: imageROM = 8'd74;
                1358: imageROM = 8'd137;
                1359: imageROM = 8'd81;
                1360: imageROM = 8'd130;
                1361: imageROM = 8'd73;
                1362: imageROM = 8'd63;
                1363: imageROM = 8'd5;
                1364: imageROM = 8'd71;
                1365: imageROM = 8'd134;
                1366: imageROM = 8'd74;
                1367: imageROM = 8'd136;
                1368: imageROM = 8'd82;
                1369: imageROM = 8'd130;
                1370: imageROM = 8'd74;
                1371: imageROM = 8'd63;
                1372: imageROM = 8'd4;
                1373: imageROM = 8'd70;
                1374: imageROM = 8'd135;
                1375: imageROM = 8'd75;
                1376: imageROM = 8'd134;
                1377: imageROM = 8'd84;
                1378: imageROM = 8'd129;
                1379: imageROM = 8'd74;
                1380: imageROM = 8'd63;
                1381: imageROM = 8'd3;
                1382: imageROM = 8'd71;
                1383: imageROM = 8'd136;
                1384: imageROM = 8'd73;
                1385: imageROM = 8'd135;
                1386: imageROM = 8'd70;
                1387: imageROM = 8'd200;
                1388: imageROM = 8'd82;
                1389: imageROM = 8'd63;
                1390: imageROM = 8'd2;
                1391: imageROM = 8'd70;
                1392: imageROM = 8'd137;
                1393: imageROM = 8'd74;
                1394: imageROM = 8'd133;
                1395: imageROM = 8'd71;
                1396: imageROM = 8'd201;
                1397: imageROM = 8'd81;
                1398: imageROM = 8'd63;
                1399: imageROM = 8'd2;
                1400: imageROM = 8'd69;
                1401: imageROM = 8'd138;
                1402: imageROM = 8'd74;
                1403: imageROM = 8'd133;
                1404: imageROM = 8'd70;
                1405: imageROM = 8'd202;
                1406: imageROM = 8'd82;
                1407: imageROM = 8'd63;
                1408: imageROM = 8'd70;
                1409: imageROM = 8'd138;
                1410: imageROM = 8'd74;
                1411: imageROM = 8'd133;
                1412: imageROM = 8'd70;
                1413: imageROM = 8'd203;
                1414: imageROM = 8'd81;
                1415: imageROM = 8'd63;
                1416: imageROM = 8'd70;
                1417: imageROM = 8'd138;
                1418: imageROM = 8'd73;
                1419: imageROM = 8'd133;
                1420: imageROM = 8'd70;
                1421: imageROM = 8'd204;
                1422: imageROM = 8'd70;
                1423: imageROM = 8'd129;
                1424: imageROM = 8'd75;
                1425: imageROM = 8'd61;
                1426: imageROM = 8'd70;
                1427: imageROM = 8'd140;
                1428: imageROM = 8'd72;
                1429: imageROM = 8'd133;
                1430: imageROM = 8'd70;
                1431: imageROM = 8'd204;
                1432: imageROM = 8'd70;
                1433: imageROM = 8'd131;
                1434: imageROM = 8'd66;
                1435: imageROM = 8'd129;
                1436: imageROM = 8'd70;
                1437: imageROM = 8'd61;
                1438: imageROM = 8'd70;
                1439: imageROM = 8'd141;
                1440: imageROM = 8'd70;
                1441: imageROM = 8'd134;
                1442: imageROM = 8'd70;
                1443: imageROM = 8'd205;
                1444: imageROM = 8'd69;
                1445: imageROM = 8'd134;
                1446: imageROM = 8'd70;
                1447: imageROM = 8'd61;
                1448: imageROM = 8'd70;
                1449: imageROM = 8'd153;
                1450: imageROM = 8'd70;
                1451: imageROM = 8'd205;
                1452: imageROM = 8'd70;
                1453: imageROM = 8'd134;
                1454: imageROM = 8'd70;
                1455: imageROM = 8'd60;
                1456: imageROM = 8'd69;
                1457: imageROM = 8'd154;
                1458: imageROM = 8'd70;
                1459: imageROM = 8'd205;
                1460: imageROM = 8'd70;
                1461: imageROM = 8'd134;
                1462: imageROM = 8'd70;
                1463: imageROM = 8'd59;
                1464: imageROM = 8'd70;
                1465: imageROM = 8'd154;
                1466: imageROM = 8'd70;
                1467: imageROM = 8'd205;
                1468: imageROM = 8'd70;
                1469: imageROM = 8'd135;
                1470: imageROM = 8'd70;
                1471: imageROM = 8'd58;
                1472: imageROM = 8'd70;
                1473: imageROM = 8'd154;
                1474: imageROM = 8'd70;
                1475: imageROM = 8'd205;
                1476: imageROM = 8'd70;
                1477: imageROM = 8'd135;
                1478: imageROM = 8'd71;
                1479: imageROM = 8'd57;
                1480: imageROM = 8'd70;
                1481: imageROM = 8'd154;
                1482: imageROM = 8'd70;
                1483: imageROM = 8'd205;
                1484: imageROM = 8'd70;
                1485: imageROM = 8'd136;
                1486: imageROM = 8'd71;
                1487: imageROM = 8'd56;
                1488: imageROM = 8'd69;
                1489: imageROM = 8'd155;
                1490: imageROM = 8'd70;
                1491: imageROM = 8'd205;
                1492: imageROM = 8'd70;
                1493: imageROM = 8'd136;
                1494: imageROM = 8'd72;
                1495: imageROM = 8'd54;
                1496: imageROM = 8'd70;
                1497: imageROM = 8'd155;
                1498: imageROM = 8'd70;
                1499: imageROM = 8'd205;
                1500: imageROM = 8'd70;
                1501: imageROM = 8'd137;
                1502: imageROM = 8'd72;
                1503: imageROM = 8'd53;
                1504: imageROM = 8'd70;
                1505: imageROM = 8'd155;
                1506: imageROM = 8'd70;
                1507: imageROM = 8'd205;
                1508: imageROM = 8'd70;
                1509: imageROM = 8'd138;
                1510: imageROM = 8'd72;
                1511: imageROM = 8'd52;
                1512: imageROM = 8'd70;
                1513: imageROM = 8'd155;
                1514: imageROM = 8'd70;
                1515: imageROM = 8'd205;
                1516: imageROM = 8'd70;
                1517: imageROM = 8'd139;
                1518: imageROM = 8'd71;
                1519: imageROM = 8'd52;
                1520: imageROM = 8'd69;
                1521: imageROM = 8'd156;
                1522: imageROM = 8'd70;
                1523: imageROM = 8'd205;
                1524: imageROM = 8'd70;
                1525: imageROM = 8'd140;
                1526: imageROM = 8'd71;
                1527: imageROM = 8'd51;
                1528: imageROM = 8'd69;
                1529: imageROM = 8'd156;
                1530: imageROM = 8'd70;
                1531: imageROM = 8'd205;
                1532: imageROM = 8'd70;
                1533: imageROM = 8'd141;
                1534: imageROM = 8'd71;
                1535: imageROM = 8'd49;
                1536: imageROM = 8'd70;
                1537: imageROM = 8'd157;
                1538: imageROM = 8'd69;
                1539: imageROM = 8'd205;
                1540: imageROM = 8'd70;
                1541: imageROM = 8'd142;
                1542: imageROM = 8'd70;
                1543: imageROM = 8'd49;
                1544: imageROM = 8'd70;
                1545: imageROM = 8'd157;
                1546: imageROM = 8'd70;
                1547: imageROM = 8'd204;
                1548: imageROM = 8'd70;
                1549: imageROM = 8'd143;
                1550: imageROM = 8'd70;
                1551: imageROM = 8'd48;
                1552: imageROM = 8'd69;
                1553: imageROM = 8'd158;
                1554: imageROM = 8'd70;
                1555: imageROM = 8'd204;
                1556: imageROM = 8'd70;
                1557: imageROM = 8'd143;
                1558: imageROM = 8'd70;
                1559: imageROM = 8'd48;
                1560: imageROM = 8'd69;
                1561: imageROM = 8'd158;
                1562: imageROM = 8'd70;
                1563: imageROM = 8'd203;
                1564: imageROM = 8'd70;
                1565: imageROM = 8'd145;
                1566: imageROM = 8'd69;
                1567: imageROM = 8'd48;
                1568: imageROM = 8'd69;
                1569: imageROM = 8'd159;
                1570: imageROM = 8'd70;
                1571: imageROM = 8'd202;
                1572: imageROM = 8'd70;
                1573: imageROM = 8'd145;
                1574: imageROM = 8'd70;
                1575: imageROM = 8'd47;
                1576: imageROM = 8'd69;
                1577: imageROM = 8'd159;
                1578: imageROM = 8'd70;
                1579: imageROM = 8'd202;
                1580: imageROM = 8'd70;
                1581: imageROM = 8'd145;
                1582: imageROM = 8'd70;
                1583: imageROM = 8'd46;
                1584: imageROM = 8'd70;
                1585: imageROM = 8'd159;
                1586: imageROM = 8'd70;
                1587: imageROM = 8'd201;
                1588: imageROM = 8'd70;
                1589: imageROM = 8'd146;
                1590: imageROM = 8'd70;
                1591: imageROM = 8'd46;
                1592: imageROM = 8'd70;
                1593: imageROM = 8'd160;
                1594: imageROM = 8'd70;
                1595: imageROM = 8'd199;
                1596: imageROM = 8'd71;
                1597: imageROM = 8'd146;
                1598: imageROM = 8'd70;
                1599: imageROM = 8'd46;
                1600: imageROM = 8'd70;
                1601: imageROM = 8'd160;
                1602: imageROM = 8'd70;
                1603: imageROM = 8'd199;
                1604: imageROM = 8'd71;
                1605: imageROM = 8'd147;
                1606: imageROM = 8'd69;
                1607: imageROM = 8'd46;
                1608: imageROM = 8'd69;
                1609: imageROM = 8'd162;
                1610: imageROM = 8'd70;
                1611: imageROM = 8'd197;
                1612: imageROM = 8'd71;
                1613: imageROM = 8'd147;
                1614: imageROM = 8'd70;
                1615: imageROM = 8'd46;
                1616: imageROM = 8'd69;
                1617: imageROM = 8'd162;
                1618: imageROM = 8'd71;
                1619: imageROM = 8'd196;
                1620: imageROM = 8'd70;
                1621: imageROM = 8'd148;
                1622: imageROM = 8'd70;
                1623: imageROM = 8'd46;
                1624: imageROM = 8'd69;
                1625: imageROM = 8'd163;
                1626: imageROM = 8'd71;
                1627: imageROM = 8'd194;
                1628: imageROM = 8'd71;
                1629: imageROM = 8'd148;
                1630: imageROM = 8'd70;
                1631: imageROM = 8'd46;
                1632: imageROM = 8'd69;
                1633: imageROM = 8'd163;
                1634: imageROM = 8'd71;
                1635: imageROM = 8'd193;
                1636: imageROM = 8'd71;
                1637: imageROM = 8'd149;
                1638: imageROM = 8'd70;
                1639: imageROM = 8'd46;
                1640: imageROM = 8'd69;
                1641: imageROM = 8'd164;
                1642: imageROM = 8'd77;
                1643: imageROM = 8'd150;
                1644: imageROM = 8'd70;
                1645: imageROM = 8'd46;
                1646: imageROM = 8'd69;
                1647: imageROM = 8'd165;
                1648: imageROM = 8'd76;
                1649: imageROM = 8'd150;
                1650: imageROM = 8'd70;
                1651: imageROM = 8'd46;
                1652: imageROM = 8'd70;
                1653: imageROM = 8'd165;
                1654: imageROM = 8'd74;
                1655: imageROM = 8'd151;
                1656: imageROM = 8'd70;
                1657: imageROM = 8'd46;
                1658: imageROM = 8'd70;
                1659: imageROM = 8'd165;
                1660: imageROM = 8'd74;
                1661: imageROM = 8'd151;
                1662: imageROM = 8'd70;
                1663: imageROM = 8'd46;
                1664: imageROM = 8'd70;
                1665: imageROM = 8'd166;
                1666: imageROM = 8'd72;
                1667: imageROM = 8'd152;
                1668: imageROM = 8'd70;
                1669: imageROM = 8'd46;
                1670: imageROM = 8'd70;
                1671: imageROM = 8'd167;
                1672: imageROM = 8'd71;
                1673: imageROM = 8'd152;
                1674: imageROM = 8'd70;
                1675: imageROM = 8'd46;
                1676: imageROM = 8'd70;
                1677: imageROM = 8'd167;
                1678: imageROM = 8'd70;
                1679: imageROM = 8'd153;
                1680: imageROM = 8'd70;
                1681: imageROM = 8'd47;
                1682: imageROM = 8'd70;
                1683: imageROM = 8'd167;
                1684: imageROM = 8'd69;
                1685: imageROM = 8'd154;
                1686: imageROM = 8'd69;
                1687: imageROM = 8'd47;
                1688: imageROM = 8'd70;
                1689: imageROM = 8'd168;
                1690: imageROM = 8'd67;
                1691: imageROM = 8'd155;
                1692: imageROM = 8'd69;
                1693: imageROM = 8'd47;
                1694: imageROM = 8'd70;
                1695: imageROM = 8'd169;
                1696: imageROM = 8'd66;
                1697: imageROM = 8'd155;
                1698: imageROM = 8'd70;
                1699: imageROM = 8'd47;
                1700: imageROM = 8'd70;
                1701: imageROM = 8'd191;
                1702: imageROM = 8'd134;
                1703: imageROM = 8'd70;
                1704: imageROM = 8'd47;
                1705: imageROM = 8'd70;
                1706: imageROM = 8'd191;
                1707: imageROM = 8'd135;
                1708: imageROM = 8'd70;
                1709: imageROM = 8'd46;
                1710: imageROM = 8'd71;
                1711: imageROM = 8'd191;
                1712: imageROM = 8'd134;
                1713: imageROM = 8'd71;
                1714: imageROM = 8'd45;
                1715: imageROM = 8'd71;
                1716: imageROM = 8'd191;
                1717: imageROM = 8'd135;
                1718: imageROM = 8'd71;
                1719: imageROM = 8'd45;
                1720: imageROM = 8'd71;
                1721: imageROM = 8'd191;
                1722: imageROM = 8'd135;
                1723: imageROM = 8'd72;
                1724: imageROM = 8'd43;
                1725: imageROM = 8'd71;
                1726: imageROM = 8'd191;
                1727: imageROM = 8'd135;
                1728: imageROM = 8'd73;
                1729: imageROM = 8'd42;
                1730: imageROM = 8'd72;
                1731: imageROM = 8'd191;
                1732: imageROM = 8'd135;
                1733: imageROM = 8'd74;
                1734: imageROM = 8'd40;
                1735: imageROM = 8'd73;
                1736: imageROM = 8'd191;
                1737: imageROM = 8'd135;
                1738: imageROM = 8'd75;
                1739: imageROM = 8'd38;
                1740: imageROM = 8'd73;
                1741: imageROM = 8'd191;
                1742: imageROM = 8'd137;
                1743: imageROM = 8'd74;
                1744: imageROM = 8'd37;
                1745: imageROM = 8'd74;
                1746: imageROM = 8'd191;
                1747: imageROM = 8'd137;
                1748: imageROM = 8'd75;
                1749: imageROM = 8'd36;
                1750: imageROM = 8'd74;
                1751: imageROM = 8'd191;
                1752: imageROM = 8'd138;
                1753: imageROM = 8'd74;
                1754: imageROM = 8'd35;
                1755: imageROM = 8'd75;
                1756: imageROM = 8'd191;
                1757: imageROM = 8'd139;
                1758: imageROM = 8'd73;
                1759: imageROM = 8'd34;
                1760: imageROM = 8'd76;
                1761: imageROM = 8'd191;
                1762: imageROM = 8'd139;
                1763: imageROM = 8'd73;
                1764: imageROM = 8'd32;
                1765: imageROM = 8'd70;
                1766: imageROM = 8'd129;
                1767: imageROM = 8'd71;
                1768: imageROM = 8'd191;
                1769: imageROM = 8'd140;
                1770: imageROM = 8'd72;
                1771: imageROM = 8'd31;
                1772: imageROM = 8'd70;
                1773: imageROM = 8'd130;
                1774: imageROM = 8'd72;
                1775: imageROM = 8'd191;
                1776: imageROM = 8'd139;
                1777: imageROM = 8'd72;
                1778: imageROM = 8'd30;
                1779: imageROM = 8'd70;
                1780: imageROM = 8'd131;
                1781: imageROM = 8'd73;
                1782: imageROM = 8'd191;
                1783: imageROM = 8'd138;
                1784: imageROM = 8'd72;
                1785: imageROM = 8'd29;
                1786: imageROM = 8'd70;
                1787: imageROM = 8'd132;
                1788: imageROM = 8'd74;
                1789: imageROM = 8'd191;
                1790: imageROM = 8'd138;
                1791: imageROM = 8'd71;
                1792: imageROM = 8'd28;
                1793: imageROM = 8'd69;
                1794: imageROM = 8'd134;
                1795: imageROM = 8'd82;
                1796: imageROM = 8'd191;
                1797: imageROM = 8'd129;
                1798: imageROM = 8'd71;
                1799: imageROM = 8'd27;
                1800: imageROM = 8'd70;
                1801: imageROM = 8'd136;
                1802: imageROM = 8'd80;
                1803: imageROM = 8'd191;
                1804: imageROM = 8'd130;
                1805: imageROM = 8'd71;
                1806: imageROM = 8'd26;
                1807: imageROM = 8'd70;
                1808: imageROM = 8'd137;
                1809: imageROM = 8'd80;
                1810: imageROM = 8'd191;
                1811: imageROM = 8'd130;
                1812: imageROM = 8'd70;
                1813: imageROM = 8'd25;
                1814: imageROM = 8'd70;
                1815: imageROM = 8'd140;
                1816: imageROM = 8'd78;
                1817: imageROM = 8'd191;
                1818: imageROM = 8'd131;
                1819: imageROM = 8'd70;
                1820: imageROM = 8'd24;
                1821: imageROM = 8'd70;
                1822: imageROM = 8'd142;
                1823: imageROM = 8'd76;
                1824: imageROM = 8'd191;
                1825: imageROM = 8'd131;
                1826: imageROM = 8'd71;
                1827: imageROM = 8'd22;
                1828: imageROM = 8'd70;
                1829: imageROM = 8'd146;
                1830: imageROM = 8'd73;
                1831: imageROM = 8'd191;
                1832: imageROM = 8'd132;
                1833: imageROM = 8'd70;
                1834: imageROM = 8'd21;
                1835: imageROM = 8'd71;
                1836: imageROM = 8'd191;
                1837: imageROM = 8'd160;
                1838: imageROM = 8'd70;
                1839: imageROM = 8'd20;
                1840: imageROM = 8'd70;
                1841: imageROM = 8'd191;
                1842: imageROM = 8'd161;
                1843: imageROM = 8'd70;
                1844: imageROM = 8'd19;
                1845: imageROM = 8'd71;
                1846: imageROM = 8'd191;
                1847: imageROM = 8'd161;
                1848: imageROM = 8'd70;
                1849: imageROM = 8'd18;
                1850: imageROM = 8'd71;
                1851: imageROM = 8'd191;
                1852: imageROM = 8'd163;
                1853: imageROM = 8'd70;
                1854: imageROM = 8'd17;
                1855: imageROM = 8'd70;
                1856: imageROM = 8'd191;
                1857: imageROM = 8'd164;
                1858: imageROM = 8'd70;
                1859: imageROM = 8'd16;
                1860: imageROM = 8'd71;
                1861: imageROM = 8'd191;
                1862: imageROM = 8'd164;
                1863: imageROM = 8'd70;
                1864: imageROM = 8'd16;
                1865: imageROM = 8'd70;
                1866: imageROM = 8'd191;
                1867: imageROM = 8'd166;
                1868: imageROM = 8'd70;
                1869: imageROM = 8'd15;
                1870: imageROM = 8'd69;
                1871: imageROM = 8'd191;
                1872: imageROM = 8'd167;
                1873: imageROM = 8'd70;
                1874: imageROM = 8'd14;
                1875: imageROM = 8'd70;
                1876: imageROM = 8'd191;
                1877: imageROM = 8'd167;
                1878: imageROM = 8'd70;
                1879: imageROM = 8'd14;
                1880: imageROM = 8'd70;
                1881: imageROM = 8'd191;
                1882: imageROM = 8'd168;
                1883: imageROM = 8'd69;
                1884: imageROM = 8'd14;
                1885: imageROM = 8'd70;
                1886: imageROM = 8'd191;
                1887: imageROM = 8'd168;
                1888: imageROM = 8'd70;
                1889: imageROM = 8'd13;
                1890: imageROM = 8'd69;
                1891: imageROM = 8'd191;
                1892: imageROM = 8'd169;
                1893: imageROM = 8'd69;
                1894: imageROM = 8'd13;
                1895: imageROM = 8'd70;
                1896: imageROM = 8'd191;
                1897: imageROM = 8'd169;
                1898: imageROM = 8'd69;
            // r04.bmp
                1899: imageROM = 8'd63;
                1900: imageROM = 8'd63;
                1901: imageROM = 8'd63;
                1902: imageROM = 8'd63;
                1903: imageROM = 8'd63;
                1904: imageROM = 8'd63;
                1905: imageROM = 8'd63;
                1906: imageROM = 8'd63;
                1907: imageROM = 8'd63;
                1908: imageROM = 8'd63;
                1909: imageROM = 8'd63;
                1910: imageROM = 8'd63;
                1911: imageROM = 8'd63;
                1912: imageROM = 8'd63;
                1913: imageROM = 8'd42;
                1914: imageROM = 8'd80;
                1915: imageROM = 8'd63;
                1916: imageROM = 8'd45;
                1917: imageROM = 8'd90;
                1918: imageROM = 8'd63;
                1919: imageROM = 8'd37;
                1920: imageROM = 8'd96;
                1921: imageROM = 8'd63;
                1922: imageROM = 8'd31;
                1923: imageROM = 8'd100;
                1924: imageROM = 8'd63;
                1925: imageROM = 8'd28;
                1926: imageROM = 8'd103;
                1927: imageROM = 8'd63;
                1928: imageROM = 8'd25;
                1929: imageROM = 8'd106;
                1930: imageROM = 8'd63;
                1931: imageROM = 8'd21;
                1932: imageROM = 8'd75;
                1933: imageROM = 8'd148;
                1934: imageROM = 8'd79;
                1935: imageROM = 8'd63;
                1936: imageROM = 8'd18;
                1937: imageROM = 8'd73;
                1938: imageROM = 8'd155;
                1939: imageROM = 8'd76;
                1940: imageROM = 8'd63;
                1941: imageROM = 8'd16;
                1942: imageROM = 8'd72;
                1943: imageROM = 8'd160;
                1944: imageROM = 8'd74;
                1945: imageROM = 8'd63;
                1946: imageROM = 8'd15;
                1947: imageROM = 8'd71;
                1948: imageROM = 8'd163;
                1949: imageROM = 8'd73;
                1950: imageROM = 8'd63;
                1951: imageROM = 8'd13;
                1952: imageROM = 8'd71;
                1953: imageROM = 8'd166;
                1954: imageROM = 8'd72;
                1955: imageROM = 8'd63;
                1956: imageROM = 8'd11;
                1957: imageROM = 8'd71;
                1958: imageROM = 8'd168;
                1959: imageROM = 8'd72;
                1960: imageROM = 8'd63;
                1961: imageROM = 8'd9;
                1962: imageROM = 8'd71;
                1963: imageROM = 8'd171;
                1964: imageROM = 8'd71;
                1965: imageROM = 8'd63;
                1966: imageROM = 8'd8;
                1967: imageROM = 8'd70;
                1968: imageROM = 8'd173;
                1969: imageROM = 8'd71;
                1970: imageROM = 8'd63;
                1971: imageROM = 8'd6;
                1972: imageROM = 8'd71;
                1973: imageROM = 8'd174;
                1974: imageROM = 8'd70;
                1975: imageROM = 8'd63;
                1976: imageROM = 8'd6;
                1977: imageROM = 8'd70;
                1978: imageROM = 8'd132;
                1979: imageROM = 8'd69;
                1980: imageROM = 8'd149;
                1981: imageROM = 8'd66;
                1982: imageROM = 8'd143;
                1983: imageROM = 8'd71;
                1984: imageROM = 8'd63;
                1985: imageROM = 8'd4;
                1986: imageROM = 8'd70;
                1987: imageROM = 8'd132;
                1988: imageROM = 8'd71;
                1989: imageROM = 8'd143;
                1990: imageROM = 8'd75;
                1991: imageROM = 8'd134;
                1992: imageROM = 8'd68;
                1993: imageROM = 8'd130;
                1994: imageROM = 8'd70;
                1995: imageROM = 8'd63;
                1996: imageROM = 8'd4;
                1997: imageROM = 8'd70;
                1998: imageROM = 8'd132;
                1999: imageROM = 8'd72;
                2000: imageROM = 8'd141;
                2001: imageROM = 8'd77;
                2002: imageROM = 8'd132;
                2003: imageROM = 8'd70;
                2004: imageROM = 8'd130;
                2005: imageROM = 8'd70;
                2006: imageROM = 8'd63;
                2007: imageROM = 8'd2;
                2008: imageROM = 8'd70;
                2009: imageROM = 8'd132;
                2010: imageROM = 8'd73;
                2011: imageROM = 8'd139;
                2012: imageROM = 8'd80;
                2013: imageROM = 8'd130;
                2014: imageROM = 8'd71;
                2015: imageROM = 8'd130;
                2016: imageROM = 8'd70;
                2017: imageROM = 8'd63;
                2018: imageROM = 8'd2;
                2019: imageROM = 8'd70;
                2020: imageROM = 8'd132;
                2021: imageROM = 8'd74;
                2022: imageROM = 8'd138;
                2023: imageROM = 8'd81;
                2024: imageROM = 8'd129;
                2025: imageROM = 8'd72;
                2026: imageROM = 8'd130;
                2027: imageROM = 8'd70;
                2028: imageROM = 8'd63;
                2029: imageROM = 8'd70;
                2030: imageROM = 8'd133;
                2031: imageROM = 8'd74;
                2032: imageROM = 8'd137;
                2033: imageROM = 8'd82;
                2034: imageROM = 8'd129;
                2035: imageROM = 8'd72;
                2036: imageROM = 8'd130;
                2037: imageROM = 8'd70;
                2038: imageROM = 8'd63;
                2039: imageROM = 8'd70;
                2040: imageROM = 8'd133;
                2041: imageROM = 8'd74;
                2042: imageROM = 8'd136;
                2043: imageROM = 8'd72;
                2044: imageROM = 8'd197;
                2045: imageROM = 8'd79;
                2046: imageROM = 8'd131;
                2047: imageROM = 8'd69;
                2048: imageROM = 8'd62;
                2049: imageROM = 8'd70;
                2050: imageROM = 8'd134;
                2051: imageROM = 8'd74;
                2052: imageROM = 8'd136;
                2053: imageROM = 8'd70;
                2054: imageROM = 8'd200;
                2055: imageROM = 8'd78;
                2056: imageROM = 8'd131;
                2057: imageROM = 8'd70;
                2058: imageROM = 8'd61;
                2059: imageROM = 8'd70;
                2060: imageROM = 8'd134;
                2061: imageROM = 8'd74;
                2062: imageROM = 8'd135;
                2063: imageROM = 8'd71;
                2064: imageROM = 8'd201;
                2065: imageROM = 8'd77;
                2066: imageROM = 8'd131;
                2067: imageROM = 8'd70;
                2068: imageROM = 8'd60;
                2069: imageROM = 8'd70;
                2070: imageROM = 8'd135;
                2071: imageROM = 8'd74;
                2072: imageROM = 8'd135;
                2073: imageROM = 8'd70;
                2074: imageROM = 8'd202;
                2075: imageROM = 8'd76;
                2076: imageROM = 8'd133;
                2077: imageROM = 8'd70;
                2078: imageROM = 8'd59;
                2079: imageROM = 8'd70;
                2080: imageROM = 8'd136;
                2081: imageROM = 8'd73;
                2082: imageROM = 8'd135;
                2083: imageROM = 8'd70;
                2084: imageROM = 8'd203;
                2085: imageROM = 8'd75;
                2086: imageROM = 8'd133;
                2087: imageROM = 8'd71;
                2088: imageROM = 8'd58;
                2089: imageROM = 8'd69;
                2090: imageROM = 8'd138;
                2091: imageROM = 8'd71;
                2092: imageROM = 8'd136;
                2093: imageROM = 8'd69;
                2094: imageROM = 8'd204;
                2095: imageROM = 8'd70;
                2096: imageROM = 8'd130;
                2097: imageROM = 8'd66;
                2098: imageROM = 8'd135;
                2099: imageROM = 8'd71;
                2100: imageROM = 8'd56;
                2101: imageROM = 8'd70;
                2102: imageROM = 8'd139;
                2103: imageROM = 8'd70;
                2104: imageROM = 8'd135;
                2105: imageROM = 8'd70;
                2106: imageROM = 8'd204;
                2107: imageROM = 8'd70;
                2108: imageROM = 8'd140;
                2109: imageROM = 8'd70;
                2110: imageROM = 8'd56;
                2111: imageROM = 8'd70;
                2112: imageROM = 8'd152;
                2113: imageROM = 8'd70;
                2114: imageROM = 8'd205;
                2115: imageROM = 8'd70;
                2116: imageROM = 8'd139;
                2117: imageROM = 8'd71;
                2118: imageROM = 8'd55;
                2119: imageROM = 8'd69;
                2120: imageROM = 8'd153;
                2121: imageROM = 8'd70;
                2122: imageROM = 8'd205;
                2123: imageROM = 8'd70;
                2124: imageROM = 8'd140;
                2125: imageROM = 8'd71;
                2126: imageROM = 8'd53;
                2127: imageROM = 8'd70;
                2128: imageROM = 8'd153;
                2129: imageROM = 8'd70;
                2130: imageROM = 8'd205;
                2131: imageROM = 8'd70;
                2132: imageROM = 8'd141;
                2133: imageROM = 8'd70;
                2134: imageROM = 8'd53;
                2135: imageROM = 8'd70;
                2136: imageROM = 8'd153;
                2137: imageROM = 8'd70;
                2138: imageROM = 8'd205;
                2139: imageROM = 8'd70;
                2140: imageROM = 8'd142;
                2141: imageROM = 8'd70;
                2142: imageROM = 8'd51;
                2143: imageROM = 8'd70;
                2144: imageROM = 8'd154;
                2145: imageROM = 8'd70;
                2146: imageROM = 8'd205;
                2147: imageROM = 8'd70;
                2148: imageROM = 8'd142;
                2149: imageROM = 8'd70;
                2150: imageROM = 8'd51;
                2151: imageROM = 8'd70;
                2152: imageROM = 8'd154;
                2153: imageROM = 8'd70;
                2154: imageROM = 8'd205;
                2155: imageROM = 8'd70;
                2156: imageROM = 8'd143;
                2157: imageROM = 8'd70;
                2158: imageROM = 8'd50;
                2159: imageROM = 8'd70;
                2160: imageROM = 8'd154;
                2161: imageROM = 8'd70;
                2162: imageROM = 8'd205;
                2163: imageROM = 8'd70;
                2164: imageROM = 8'd143;
                2165: imageROM = 8'd70;
                2166: imageROM = 8'd49;
                2167: imageROM = 8'd70;
                2168: imageROM = 8'd155;
                2169: imageROM = 8'd70;
                2170: imageROM = 8'd205;
                2171: imageROM = 8'd70;
                2172: imageROM = 8'd144;
                2173: imageROM = 8'd69;
                2174: imageROM = 8'd49;
                2175: imageROM = 8'd70;
                2176: imageROM = 8'd155;
                2177: imageROM = 8'd70;
                2178: imageROM = 8'd205;
                2179: imageROM = 8'd70;
                2180: imageROM = 8'd144;
                2181: imageROM = 8'd70;
                2182: imageROM = 8'd48;
                2183: imageROM = 8'd70;
                2184: imageROM = 8'd155;
                2185: imageROM = 8'd70;
                2186: imageROM = 8'd205;
                2187: imageROM = 8'd70;
                2188: imageROM = 8'd144;
                2189: imageROM = 8'd70;
                2190: imageROM = 8'd48;
                2191: imageROM = 8'd70;
                2192: imageROM = 8'd155;
                2193: imageROM = 8'd70;
                2194: imageROM = 8'd205;
                2195: imageROM = 8'd70;
                2196: imageROM = 8'd144;
                2197: imageROM = 8'd70;
                2198: imageROM = 8'd48;
                2199: imageROM = 8'd69;
                2200: imageROM = 8'd157;
                2201: imageROM = 8'd69;
                2202: imageROM = 8'd205;
                2203: imageROM = 8'd70;
                2204: imageROM = 8'd145;
                2205: imageROM = 8'd69;
                2206: imageROM = 8'd48;
                2207: imageROM = 8'd69;
                2208: imageROM = 8'd157;
                2209: imageROM = 8'd70;
                2210: imageROM = 8'd204;
                2211: imageROM = 8'd70;
                2212: imageROM = 8'd145;
                2213: imageROM = 8'd69;
                2214: imageROM = 8'd47;
                2215: imageROM = 8'd70;
                2216: imageROM = 8'd157;
                2217: imageROM = 8'd70;
                2218: imageROM = 8'd204;
                2219: imageROM = 8'd70;
                2220: imageROM = 8'd145;
                2221: imageROM = 8'd69;
                2222: imageROM = 8'd47;
                2223: imageROM = 8'd70;
                2224: imageROM = 8'd157;
                2225: imageROM = 8'd70;
                2226: imageROM = 8'd204;
                2227: imageROM = 8'd69;
                2228: imageROM = 8'd146;
                2229: imageROM = 8'd69;
                2230: imageROM = 8'd47;
                2231: imageROM = 8'd70;
                2232: imageROM = 8'd158;
                2233: imageROM = 8'd70;
                2234: imageROM = 8'd202;
                2235: imageROM = 8'd70;
                2236: imageROM = 8'd146;
                2237: imageROM = 8'd69;
                2238: imageROM = 8'd47;
                2239: imageROM = 8'd70;
                2240: imageROM = 8'd158;
                2241: imageROM = 8'd70;
                2242: imageROM = 8'd202;
                2243: imageROM = 8'd70;
                2244: imageROM = 8'd146;
                2245: imageROM = 8'd69;
                2246: imageROM = 8'd47;
                2247: imageROM = 8'd70;
                2248: imageROM = 8'd158;
                2249: imageROM = 8'd70;
                2250: imageROM = 8'd202;
                2251: imageROM = 8'd70;
                2252: imageROM = 8'd146;
                2253: imageROM = 8'd69;
                2254: imageROM = 8'd47;
                2255: imageROM = 8'd70;
                2256: imageROM = 8'd159;
                2257: imageROM = 8'd70;
                2258: imageROM = 8'd200;
                2259: imageROM = 8'd70;
                2260: imageROM = 8'd147;
                2261: imageROM = 8'd69;
                2262: imageROM = 8'd47;
                2263: imageROM = 8'd70;
                2264: imageROM = 8'd159;
                2265: imageROM = 8'd70;
                2266: imageROM = 8'd199;
                2267: imageROM = 8'd71;
                2268: imageROM = 8'd147;
                2269: imageROM = 8'd69;
                2270: imageROM = 8'd47;
                2271: imageROM = 8'd70;
                2272: imageROM = 8'd160;
                2273: imageROM = 8'd70;
                2274: imageROM = 8'd198;
                2275: imageROM = 8'd70;
                2276: imageROM = 8'd147;
                2277: imageROM = 8'd70;
                2278: imageROM = 8'd47;
                2279: imageROM = 8'd70;
                2280: imageROM = 8'd160;
                2281: imageROM = 8'd71;
                2282: imageROM = 8'd196;
                2283: imageROM = 8'd71;
                2284: imageROM = 8'd147;
                2285: imageROM = 8'd70;
                2286: imageROM = 8'd47;
                2287: imageROM = 8'd70;
                2288: imageROM = 8'd161;
                2289: imageROM = 8'd70;
                2290: imageROM = 8'd195;
                2291: imageROM = 8'd71;
                2292: imageROM = 8'd148;
                2293: imageROM = 8'd70;
                2294: imageROM = 8'd47;
                2295: imageROM = 8'd70;
                2296: imageROM = 8'd161;
                2297: imageROM = 8'd71;
                2298: imageROM = 8'd194;
                2299: imageROM = 8'd70;
                2300: imageROM = 8'd149;
                2301: imageROM = 8'd69;
                2302: imageROM = 8'd48;
                2303: imageROM = 8'd70;
                2304: imageROM = 8'd162;
                2305: imageROM = 8'd71;
                2306: imageROM = 8'd193;
                2307: imageROM = 8'd70;
                2308: imageROM = 8'd149;
                2309: imageROM = 8'd69;
                2310: imageROM = 8'd48;
                2311: imageROM = 8'd70;
                2312: imageROM = 8'd163;
                2313: imageROM = 8'd76;
                2314: imageROM = 8'd150;
                2315: imageROM = 8'd69;
                2316: imageROM = 8'd48;
                2317: imageROM = 8'd70;
                2318: imageROM = 8'd164;
                2319: imageROM = 8'd75;
                2320: imageROM = 8'd150;
                2321: imageROM = 8'd69;
                2322: imageROM = 8'd48;
                2323: imageROM = 8'd70;
                2324: imageROM = 8'd164;
                2325: imageROM = 8'd74;
                2326: imageROM = 8'd151;
                2327: imageROM = 8'd69;
                2328: imageROM = 8'd49;
                2329: imageROM = 8'd70;
                2330: imageROM = 8'd164;
                2331: imageROM = 8'd72;
                2332: imageROM = 8'd152;
                2333: imageROM = 8'd69;
                2334: imageROM = 8'd49;
                2335: imageROM = 8'd70;
                2336: imageROM = 8'd165;
                2337: imageROM = 8'd71;
                2338: imageROM = 8'd152;
                2339: imageROM = 8'd70;
                2340: imageROM = 8'd48;
                2341: imageROM = 8'd70;
                2342: imageROM = 8'd165;
                2343: imageROM = 8'd70;
                2344: imageROM = 8'd153;
                2345: imageROM = 8'd70;
                2346: imageROM = 8'd48;
                2347: imageROM = 8'd70;
                2348: imageROM = 8'd166;
                2349: imageROM = 8'd69;
                2350: imageROM = 8'd154;
                2351: imageROM = 8'd69;
                2352: imageROM = 8'd48;
                2353: imageROM = 8'd71;
                2354: imageROM = 8'd166;
                2355: imageROM = 8'd67;
                2356: imageROM = 8'd155;
                2357: imageROM = 8'd70;
                2358: imageROM = 8'd48;
                2359: imageROM = 8'd70;
                2360: imageROM = 8'd166;
                2361: imageROM = 8'd67;
                2362: imageROM = 8'd155;
                2363: imageROM = 8'd71;
                2364: imageROM = 8'd47;
                2365: imageROM = 8'd70;
                2366: imageROM = 8'd167;
                2367: imageROM = 8'd66;
                2368: imageROM = 8'd156;
                2369: imageROM = 8'd70;
                2370: imageROM = 8'd48;
                2371: imageROM = 8'd70;
                2372: imageROM = 8'd191;
                2373: imageROM = 8'd134;
                2374: imageROM = 8'd70;
                2375: imageROM = 8'd47;
                2376: imageROM = 8'd70;
                2377: imageROM = 8'd191;
                2378: imageROM = 8'd134;
                2379: imageROM = 8'd71;
                2380: imageROM = 8'd47;
                2381: imageROM = 8'd70;
                2382: imageROM = 8'd191;
                2383: imageROM = 8'd134;
                2384: imageROM = 8'd71;
                2385: imageROM = 8'd46;
                2386: imageROM = 8'd71;
                2387: imageROM = 8'd191;
                2388: imageROM = 8'd133;
                2389: imageROM = 8'd72;
                2390: imageROM = 8'd46;
                2391: imageROM = 8'd70;
                2392: imageROM = 8'd191;
                2393: imageROM = 8'd134;
                2394: imageROM = 8'd72;
                2395: imageROM = 8'd45;
                2396: imageROM = 8'd71;
                2397: imageROM = 8'd191;
                2398: imageROM = 8'd134;
                2399: imageROM = 8'd72;
                2400: imageROM = 8'd45;
                2401: imageROM = 8'd71;
                2402: imageROM = 8'd191;
                2403: imageROM = 8'd134;
                2404: imageROM = 8'd72;
                2405: imageROM = 8'd44;
                2406: imageROM = 8'd71;
                2407: imageROM = 8'd191;
                2408: imageROM = 8'd135;
                2409: imageROM = 8'd73;
                2410: imageROM = 8'd43;
                2411: imageROM = 8'd71;
                2412: imageROM = 8'd191;
                2413: imageROM = 8'd135;
                2414: imageROM = 8'd73;
                2415: imageROM = 8'd42;
                2416: imageROM = 8'd72;
                2417: imageROM = 8'd191;
                2418: imageROM = 8'd135;
                2419: imageROM = 8'd74;
                2420: imageROM = 8'd40;
                2421: imageROM = 8'd73;
                2422: imageROM = 8'd191;
                2423: imageROM = 8'd135;
                2424: imageROM = 8'd75;
                2425: imageROM = 8'd38;
                2426: imageROM = 8'd74;
                2427: imageROM = 8'd191;
                2428: imageROM = 8'd136;
                2429: imageROM = 8'd75;
                2430: imageROM = 8'd36;
                2431: imageROM = 8'd76;
                2432: imageROM = 8'd191;
                2433: imageROM = 8'd135;
                2434: imageROM = 8'd77;
                2435: imageROM = 8'd33;
                2436: imageROM = 8'd77;
                2437: imageROM = 8'd191;
                2438: imageROM = 8'd136;
                2439: imageROM = 8'd77;
                2440: imageROM = 8'd31;
                2441: imageROM = 8'd79;
                2442: imageROM = 8'd191;
                2443: imageROM = 8'd136;
                2444: imageROM = 8'd77;
                2445: imageROM = 8'd29;
                2446: imageROM = 8'd69;
                2447: imageROM = 8'd131;
                2448: imageROM = 8'd72;
                2449: imageROM = 8'd191;
                2450: imageROM = 8'd137;
                2451: imageROM = 8'd77;
                2452: imageROM = 8'd27;
                2453: imageROM = 8'd69;
                2454: imageROM = 8'd132;
                2455: imageROM = 8'd73;
                2456: imageROM = 8'd191;
                2457: imageROM = 8'd137;
                2458: imageROM = 8'd77;
                2459: imageROM = 8'd25;
                2460: imageROM = 8'd69;
                2461: imageROM = 8'd133;
                2462: imageROM = 8'd75;
                2463: imageROM = 8'd191;
                2464: imageROM = 8'd137;
                2465: imageROM = 8'd75;
                2466: imageROM = 8'd24;
                2467: imageROM = 8'd69;
                2468: imageROM = 8'd134;
                2469: imageROM = 8'd82;
                2470: imageROM = 8'd191;
                2471: imageROM = 8'd131;
                2472: imageROM = 8'd75;
                2473: imageROM = 8'd21;
                2474: imageROM = 8'd70;
                2475: imageROM = 8'd136;
                2476: imageROM = 8'd80;
                2477: imageROM = 8'd191;
                2478: imageROM = 8'd133;
                2479: imageROM = 8'd74;
                2480: imageROM = 8'd20;
                2481: imageROM = 8'd70;
                2482: imageROM = 8'd138;
                2483: imageROM = 8'd79;
                2484: imageROM = 8'd191;
                2485: imageROM = 8'd134;
                2486: imageROM = 8'd73;
                2487: imageROM = 8'd19;
                2488: imageROM = 8'd70;
                2489: imageROM = 8'd140;
                2490: imageROM = 8'd77;
                2491: imageROM = 8'd191;
                2492: imageROM = 8'd136;
                2493: imageROM = 8'd72;
                2494: imageROM = 8'd18;
                2495: imageROM = 8'd70;
                2496: imageROM = 8'd143;
                2497: imageROM = 8'd74;
                2498: imageROM = 8'd191;
                2499: imageROM = 8'd137;
                2500: imageROM = 8'd71;
                2501: imageROM = 8'd18;
                2502: imageROM = 8'd69;
                2503: imageROM = 8'd149;
                2504: imageROM = 8'd67;
                2505: imageROM = 8'd191;
                2506: imageROM = 8'd140;
                2507: imageROM = 8'd71;
                2508: imageROM = 8'd17;
                2509: imageROM = 8'd69;
                2510: imageROM = 8'd191;
                2511: imageROM = 8'd165;
                2512: imageROM = 8'd71;
                2513: imageROM = 8'd16;
                2514: imageROM = 8'd69;
                2515: imageROM = 8'd191;
                2516: imageROM = 8'd166;
                2517: imageROM = 8'd70;
                2518: imageROM = 8'd16;
                2519: imageROM = 8'd69;
                2520: imageROM = 8'd191;
                2521: imageROM = 8'd167;
                2522: imageROM = 8'd70;
                2523: imageROM = 8'd15;
                2524: imageROM = 8'd69;
                2525: imageROM = 8'd191;
                2526: imageROM = 8'd167;
                2527: imageROM = 8'd71;
                2528: imageROM = 8'd14;
                2529: imageROM = 8'd69;
                2530: imageROM = 8'd191;
                2531: imageROM = 8'd168;
                2532: imageROM = 8'd70;
            // r05.bmp
                2533: imageROM = 8'd63;
                2534: imageROM = 8'd63;
                2535: imageROM = 8'd63;
                2536: imageROM = 8'd63;
                2537: imageROM = 8'd63;
                2538: imageROM = 8'd63;
                2539: imageROM = 8'd63;
                2540: imageROM = 8'd63;
                2541: imageROM = 8'd63;
                2542: imageROM = 8'd63;
                2543: imageROM = 8'd63;
                2544: imageROM = 8'd63;
                2545: imageROM = 8'd63;
                2546: imageROM = 8'd63;
                2547: imageROM = 8'd48;
                2548: imageROM = 8'd78;
                2549: imageROM = 8'd63;
                2550: imageROM = 8'd47;
                2551: imageROM = 8'd88;
                2552: imageROM = 8'd63;
                2553: imageROM = 8'd38;
                2554: imageROM = 8'd94;
                2555: imageROM = 8'd63;
                2556: imageROM = 8'd33;
                2557: imageROM = 8'd98;
                2558: imageROM = 8'd63;
                2559: imageROM = 8'd30;
                2560: imageROM = 8'd101;
                2561: imageROM = 8'd63;
                2562: imageROM = 8'd26;
                2563: imageROM = 8'd105;
                2564: imageROM = 8'd63;
                2565: imageROM = 8'd23;
                2566: imageROM = 8'd75;
                2567: imageROM = 8'd146;
                2568: imageROM = 8'd79;
                2569: imageROM = 8'd63;
                2570: imageROM = 8'd20;
                2571: imageROM = 8'd74;
                2572: imageROM = 8'd152;
                2573: imageROM = 8'd76;
                2574: imageROM = 8'd63;
                2575: imageROM = 8'd17;
                2576: imageROM = 8'd74;
                2577: imageROM = 8'd157;
                2578: imageROM = 8'd74;
                2579: imageROM = 8'd63;
                2580: imageROM = 8'd15;
                2581: imageROM = 8'd73;
                2582: imageROM = 8'd161;
                2583: imageROM = 8'd73;
                2584: imageROM = 8'd63;
                2585: imageROM = 8'd13;
                2586: imageROM = 8'd72;
                2587: imageROM = 8'd165;
                2588: imageROM = 8'd72;
                2589: imageROM = 8'd63;
                2590: imageROM = 8'd11;
                2591: imageROM = 8'd72;
                2592: imageROM = 8'd167;
                2593: imageROM = 8'd72;
                2594: imageROM = 8'd63;
                2595: imageROM = 8'd9;
                2596: imageROM = 8'd72;
                2597: imageROM = 8'd170;
                2598: imageROM = 8'd71;
                2599: imageROM = 8'd63;
                2600: imageROM = 8'd8;
                2601: imageROM = 8'd71;
                2602: imageROM = 8'd172;
                2603: imageROM = 8'd70;
                2604: imageROM = 8'd63;
                2605: imageROM = 8'd7;
                2606: imageROM = 8'd71;
                2607: imageROM = 8'd173;
                2608: imageROM = 8'd71;
                2609: imageROM = 8'd63;
                2610: imageROM = 8'd5;
                2611: imageROM = 8'd71;
                2612: imageROM = 8'd175;
                2613: imageROM = 8'd70;
                2614: imageROM = 8'd63;
                2615: imageROM = 8'd4;
                2616: imageROM = 8'd71;
                2617: imageROM = 8'd177;
                2618: imageROM = 8'd70;
                2619: imageROM = 8'd63;
                2620: imageROM = 8'd2;
                2621: imageROM = 8'd71;
                2622: imageROM = 8'd178;
                2623: imageROM = 8'd70;
                2624: imageROM = 8'd63;
                2625: imageROM = 8'd2;
                2626: imageROM = 8'd70;
                2627: imageROM = 8'd180;
                2628: imageROM = 8'd70;
                2629: imageROM = 8'd63;
                2630: imageROM = 8'd70;
                2631: imageROM = 8'd136;
                2632: imageROM = 8'd70;
                2633: imageROM = 8'd142;
                2634: imageROM = 8'd71;
                2635: imageROM = 8'd141;
                2636: imageROM = 8'd65;
                2637: imageROM = 8'd132;
                2638: imageROM = 8'd70;
                2639: imageROM = 8'd62;
                2640: imageROM = 8'd71;
                2641: imageROM = 8'd135;
                2642: imageROM = 8'd72;
                2643: imageROM = 8'd139;
                2644: imageROM = 8'd75;
                2645: imageROM = 8'd137;
                2646: imageROM = 8'd69;
                2647: imageROM = 8'd130;
                2648: imageROM = 8'd70;
                2649: imageROM = 8'd61;
                2650: imageROM = 8'd71;
                2651: imageROM = 8'd136;
                2652: imageROM = 8'd73;
                2653: imageROM = 8'd137;
                2654: imageROM = 8'd78;
                2655: imageROM = 8'd134;
                2656: imageROM = 8'd71;
                2657: imageROM = 8'd130;
                2658: imageROM = 8'd70;
                2659: imageROM = 8'd60;
                2660: imageROM = 8'd70;
                2661: imageROM = 8'd137;
                2662: imageROM = 8'd73;
                2663: imageROM = 8'd136;
                2664: imageROM = 8'd80;
                2665: imageROM = 8'd133;
                2666: imageROM = 8'd71;
                2667: imageROM = 8'd130;
                2668: imageROM = 8'd70;
                2669: imageROM = 8'd59;
                2670: imageROM = 8'd71;
                2671: imageROM = 8'd137;
                2672: imageROM = 8'd74;
                2673: imageROM = 8'd134;
                2674: imageROM = 8'd82;
                2675: imageROM = 8'd132;
                2676: imageROM = 8'd72;
                2677: imageROM = 8'd130;
                2678: imageROM = 8'd70;
                2679: imageROM = 8'd58;
                2680: imageROM = 8'd70;
                2681: imageROM = 8'd138;
                2682: imageROM = 8'd74;
                2683: imageROM = 8'd133;
                2684: imageROM = 8'd83;
                2685: imageROM = 8'd132;
                2686: imageROM = 8'd72;
                2687: imageROM = 8'd130;
                2688: imageROM = 8'd71;
                2689: imageROM = 8'd56;
                2690: imageROM = 8'd71;
                2691: imageROM = 8'd138;
                2692: imageROM = 8'd74;
                2693: imageROM = 8'd133;
                2694: imageROM = 8'd71;
                2695: imageROM = 8'd198;
                2696: imageROM = 8'd71;
                2697: imageROM = 8'd131;
                2698: imageROM = 8'd72;
                2699: imageROM = 8'd131;
                2700: imageROM = 8'd71;
                2701: imageROM = 8'd55;
                2702: imageROM = 8'd70;
                2703: imageROM = 8'd139;
                2704: imageROM = 8'd74;
                2705: imageROM = 8'd132;
                2706: imageROM = 8'd71;
                2707: imageROM = 8'd200;
                2708: imageROM = 8'd70;
                2709: imageROM = 8'd131;
                2710: imageROM = 8'd72;
                2711: imageROM = 8'd132;
                2712: imageROM = 8'd70;
                2713: imageROM = 8'd54;
                2714: imageROM = 8'd70;
                2715: imageROM = 8'd140;
                2716: imageROM = 8'd74;
                2717: imageROM = 8'd132;
                2718: imageROM = 8'd70;
                2719: imageROM = 8'd202;
                2720: imageROM = 8'd70;
                2721: imageROM = 8'd130;
                2722: imageROM = 8'd72;
                2723: imageROM = 8'd132;
                2724: imageROM = 8'd71;
                2725: imageROM = 8'd53;
                2726: imageROM = 8'd70;
                2727: imageROM = 8'd140;
                2728: imageROM = 8'd74;
                2729: imageROM = 8'd131;
                2730: imageROM = 8'd70;
                2731: imageROM = 8'd203;
                2732: imageROM = 8'd70;
                2733: imageROM = 8'd131;
                2734: imageROM = 8'd70;
                2735: imageROM = 8'd134;
                2736: imageROM = 8'd71;
                2737: imageROM = 8'd51;
                2738: imageROM = 8'd70;
                2739: imageROM = 8'd142;
                2740: imageROM = 8'd72;
                2741: imageROM = 8'd132;
                2742: imageROM = 8'd70;
                2743: imageROM = 8'd204;
                2744: imageROM = 8'd69;
                2745: imageROM = 8'd132;
                2746: imageROM = 8'd69;
                2747: imageROM = 8'd135;
                2748: imageROM = 8'd71;
                2749: imageROM = 8'd50;
                2750: imageROM = 8'd70;
                2751: imageROM = 8'd142;
                2752: imageROM = 8'd72;
                2753: imageROM = 8'd132;
                2754: imageROM = 8'd70;
                2755: imageROM = 8'd204;
                2756: imageROM = 8'd70;
                2757: imageROM = 8'd144;
                2758: imageROM = 8'd70;
                2759: imageROM = 8'd49;
                2760: imageROM = 8'd70;
                2761: imageROM = 8'd145;
                2762: imageROM = 8'd69;
                2763: imageROM = 8'd133;
                2764: imageROM = 8'd70;
                2765: imageROM = 8'd204;
                2766: imageROM = 8'd70;
                2767: imageROM = 8'd144;
                2768: imageROM = 8'd71;
                2769: imageROM = 8'd48;
                2770: imageROM = 8'd70;
                2771: imageROM = 8'd155;
                2772: imageROM = 8'd69;
                2773: imageROM = 8'd205;
                2774: imageROM = 8'd70;
                2775: imageROM = 8'd145;
                2776: imageROM = 8'd70;
                2777: imageROM = 8'd48;
                2778: imageROM = 8'd70;
                2779: imageROM = 8'd155;
                2780: imageROM = 8'd69;
                2781: imageROM = 8'd206;
                2782: imageROM = 8'd69;
                2783: imageROM = 8'd146;
                2784: imageROM = 8'd70;
                2785: imageROM = 8'd46;
                2786: imageROM = 8'd70;
                2787: imageROM = 8'd155;
                2788: imageROM = 8'd70;
                2789: imageROM = 8'd206;
                2790: imageROM = 8'd70;
                2791: imageROM = 8'd145;
                2792: imageROM = 8'd70;
                2793: imageROM = 8'd46;
                2794: imageROM = 8'd70;
                2795: imageROM = 8'd155;
                2796: imageROM = 8'd70;
                2797: imageROM = 8'd206;
                2798: imageROM = 8'd70;
                2799: imageROM = 8'd145;
                2800: imageROM = 8'd70;
                2801: imageROM = 8'd46;
                2802: imageROM = 8'd70;
                2803: imageROM = 8'd155;
                2804: imageROM = 8'd70;
                2805: imageROM = 8'd206;
                2806: imageROM = 8'd70;
                2807: imageROM = 8'd146;
                2808: imageROM = 8'd70;
                2809: imageROM = 8'd45;
                2810: imageROM = 8'd70;
                2811: imageROM = 8'd155;
                2812: imageROM = 8'd70;
                2813: imageROM = 8'd206;
                2814: imageROM = 8'd70;
                2815: imageROM = 8'd146;
                2816: imageROM = 8'd70;
                2817: imageROM = 8'd45;
                2818: imageROM = 8'd69;
                2819: imageROM = 8'd157;
                2820: imageROM = 8'd69;
                2821: imageROM = 8'd206;
                2822: imageROM = 8'd70;
                2823: imageROM = 8'd146;
                2824: imageROM = 8'd70;
                2825: imageROM = 8'd44;
                2826: imageROM = 8'd70;
                2827: imageROM = 8'd157;
                2828: imageROM = 8'd69;
                2829: imageROM = 8'd206;
                2830: imageROM = 8'd70;
                2831: imageROM = 8'd147;
                2832: imageROM = 8'd69;
                2833: imageROM = 8'd44;
                2834: imageROM = 8'd70;
                2835: imageROM = 8'd157;
                2836: imageROM = 8'd69;
                2837: imageROM = 8'd206;
                2838: imageROM = 8'd70;
                2839: imageROM = 8'd147;
                2840: imageROM = 8'd69;
                2841: imageROM = 8'd44;
                2842: imageROM = 8'd70;
                2843: imageROM = 8'd157;
                2844: imageROM = 8'd70;
                2845: imageROM = 8'd205;
                2846: imageROM = 8'd70;
                2847: imageROM = 8'd147;
                2848: imageROM = 8'd69;
                2849: imageROM = 8'd44;
                2850: imageROM = 8'd70;
                2851: imageROM = 8'd157;
                2852: imageROM = 8'd70;
                2853: imageROM = 8'd205;
                2854: imageROM = 8'd70;
                2855: imageROM = 8'd147;
                2856: imageROM = 8'd70;
                2857: imageROM = 8'd43;
                2858: imageROM = 8'd69;
                2859: imageROM = 8'd158;
                2860: imageROM = 8'd70;
                2861: imageROM = 8'd205;
                2862: imageROM = 8'd70;
                2863: imageROM = 8'd147;
                2864: imageROM = 8'd70;
                2865: imageROM = 8'd43;
                2866: imageROM = 8'd69;
                2867: imageROM = 8'd158;
                2868: imageROM = 8'd70;
                2869: imageROM = 8'd205;
                2870: imageROM = 8'd69;
                2871: imageROM = 8'd148;
                2872: imageROM = 8'd70;
                2873: imageROM = 8'd43;
                2874: imageROM = 8'd69;
                2875: imageROM = 8'd159;
                2876: imageROM = 8'd70;
                2877: imageROM = 8'd203;
                2878: imageROM = 8'd70;
                2879: imageROM = 8'd148;
                2880: imageROM = 8'd69;
                2881: imageROM = 8'd44;
                2882: imageROM = 8'd69;
                2883: imageROM = 8'd159;
                2884: imageROM = 8'd70;
                2885: imageROM = 8'd203;
                2886: imageROM = 8'd70;
                2887: imageROM = 8'd148;
                2888: imageROM = 8'd69;
                2889: imageROM = 8'd44;
                2890: imageROM = 8'd69;
                2891: imageROM = 8'd159;
                2892: imageROM = 8'd70;
                2893: imageROM = 8'd203;
                2894: imageROM = 8'd70;
                2895: imageROM = 8'd148;
                2896: imageROM = 8'd69;
                2897: imageROM = 8'd44;
                2898: imageROM = 8'd69;
                2899: imageROM = 8'd159;
                2900: imageROM = 8'd71;
                2901: imageROM = 8'd202;
                2902: imageROM = 8'd69;
                2903: imageROM = 8'd148;
                2904: imageROM = 8'd70;
                2905: imageROM = 8'd44;
                2906: imageROM = 8'd69;
                2907: imageROM = 8'd160;
                2908: imageROM = 8'd70;
                2909: imageROM = 8'd201;
                2910: imageROM = 8'd70;
                2911: imageROM = 8'd148;
                2912: imageROM = 8'd70;
                2913: imageROM = 8'd44;
                2914: imageROM = 8'd69;
                2915: imageROM = 8'd160;
                2916: imageROM = 8'd70;
                2917: imageROM = 8'd200;
                2918: imageROM = 8'd71;
                2919: imageROM = 8'd148;
                2920: imageROM = 8'd70;
                2921: imageROM = 8'd44;
                2922: imageROM = 8'd70;
                2923: imageROM = 8'd160;
                2924: imageROM = 8'd70;
                2925: imageROM = 8'd199;
                2926: imageROM = 8'd70;
                2927: imageROM = 8'd149;
                2928: imageROM = 8'd70;
                2929: imageROM = 8'd44;
                2930: imageROM = 8'd70;
                2931: imageROM = 8'd160;
                2932: imageROM = 8'd71;
                2933: imageROM = 8'd197;
                2934: imageROM = 8'd71;
                2935: imageROM = 8'd149;
                2936: imageROM = 8'd69;
                2937: imageROM = 8'd45;
                2938: imageROM = 8'd70;
                2939: imageROM = 8'd160;
                2940: imageROM = 8'd71;
                2941: imageROM = 8'd196;
                2942: imageROM = 8'd71;
                2943: imageROM = 8'd149;
                2944: imageROM = 8'd70;
                2945: imageROM = 8'd45;
                2946: imageROM = 8'd70;
                2947: imageROM = 8'd161;
                2948: imageROM = 8'd71;
                2949: imageROM = 8'd195;
                2950: imageROM = 8'd70;
                2951: imageROM = 8'd150;
                2952: imageROM = 8'd70;
                2953: imageROM = 8'd45;
                2954: imageROM = 8'd70;
                2955: imageROM = 8'd162;
                2956: imageROM = 8'd71;
                2957: imageROM = 8'd193;
                2958: imageROM = 8'd71;
                2959: imageROM = 8'd150;
                2960: imageROM = 8'd70;
                2961: imageROM = 8'd46;
                2962: imageROM = 8'd69;
                2963: imageROM = 8'd163;
                2964: imageROM = 8'd70;
                2965: imageROM = 8'd193;
                2966: imageROM = 8'd70;
                2967: imageROM = 8'd152;
                2968: imageROM = 8'd69;
                2969: imageROM = 8'd46;
                2970: imageROM = 8'd69;
                2971: imageROM = 8'd163;
                2972: imageROM = 8'd77;
                2973: imageROM = 8'd152;
                2974: imageROM = 8'd70;
                2975: imageROM = 8'd45;
                2976: imageROM = 8'd70;
                2977: imageROM = 8'd163;
                2978: imageROM = 8'd75;
                2979: imageROM = 8'd153;
                2980: imageROM = 8'd70;
                2981: imageROM = 8'd45;
                2982: imageROM = 8'd70;
                2983: imageROM = 8'd164;
                2984: imageROM = 8'd74;
                2985: imageROM = 8'd154;
                2986: imageROM = 8'd70;
                2987: imageROM = 8'd44;
                2988: imageROM = 8'd70;
                2989: imageROM = 8'd165;
                2990: imageROM = 8'd72;
                2991: imageROM = 8'd155;
                2992: imageROM = 8'd70;
                2993: imageROM = 8'd44;
                2994: imageROM = 8'd70;
                2995: imageROM = 8'd165;
                2996: imageROM = 8'd71;
                2997: imageROM = 8'd157;
                2998: imageROM = 8'd70;
                2999: imageROM = 8'd43;
                3000: imageROM = 8'd71;
                3001: imageROM = 8'd165;
                3002: imageROM = 8'd70;
                3003: imageROM = 8'd157;
                3004: imageROM = 8'd71;
                3005: imageROM = 8'd43;
                3006: imageROM = 8'd70;
                3007: imageROM = 8'd166;
                3008: imageROM = 8'd68;
                3009: imageROM = 8'd159;
                3010: imageROM = 8'd70;
                3011: imageROM = 8'd43;
                3012: imageROM = 8'd70;
                3013: imageROM = 8'd166;
                3014: imageROM = 8'd68;
                3015: imageROM = 8'd159;
                3016: imageROM = 8'd71;
                3017: imageROM = 8'd42;
                3018: imageROM = 8'd71;
                3019: imageROM = 8'd166;
                3020: imageROM = 8'd67;
                3021: imageROM = 8'd160;
                3022: imageROM = 8'd71;
                3023: imageROM = 8'd41;
                3024: imageROM = 8'd71;
                3025: imageROM = 8'd167;
                3026: imageROM = 8'd65;
                3027: imageROM = 8'd162;
                3028: imageROM = 8'd71;
                3029: imageROM = 8'd40;
                3030: imageROM = 8'd72;
                3031: imageROM = 8'd191;
                3032: imageROM = 8'd139;
                3033: imageROM = 8'd71;
                3034: imageROM = 8'd40;
                3035: imageROM = 8'd72;
                3036: imageROM = 8'd191;
                3037: imageROM = 8'd139;
                3038: imageROM = 8'd72;
                3039: imageROM = 8'd38;
                3040: imageROM = 8'd72;
                3041: imageROM = 8'd191;
                3042: imageROM = 8'd140;
                3043: imageROM = 8'd72;
                3044: imageROM = 8'd37;
                3045: imageROM = 8'd73;
                3046: imageROM = 8'd191;
                3047: imageROM = 8'd140;
                3048: imageROM = 8'd73;
                3049: imageROM = 8'd35;
                3050: imageROM = 8'd74;
                3051: imageROM = 8'd191;
                3052: imageROM = 8'd140;
                3053: imageROM = 8'd73;
                3054: imageROM = 8'd34;
                3055: imageROM = 8'd75;
                3056: imageROM = 8'd191;
                3057: imageROM = 8'd140;
                3058: imageROM = 8'd74;
                3059: imageROM = 8'd32;
                3060: imageROM = 8'd76;
                3061: imageROM = 8'd191;
                3062: imageROM = 8'd140;
                3063: imageROM = 8'd76;
                3064: imageROM = 8'd29;
                3065: imageROM = 8'd77;
                3066: imageROM = 8'd191;
                3067: imageROM = 8'd141;
                3068: imageROM = 8'd76;
                3069: imageROM = 8'd27;
                3070: imageROM = 8'd78;
                3071: imageROM = 8'd191;
                3072: imageROM = 8'd141;
                3073: imageROM = 8'd77;
                3074: imageROM = 8'd25;
                3075: imageROM = 8'd70;
                3076: imageROM = 8'd129;
                3077: imageROM = 8'd72;
                3078: imageROM = 8'd191;
                3079: imageROM = 8'd142;
                3080: imageROM = 8'd78;
                3081: imageROM = 8'd23;
                3082: imageROM = 8'd69;
                3083: imageROM = 8'd130;
                3084: imageROM = 8'd73;
                3085: imageROM = 8'd191;
                3086: imageROM = 8'd142;
                3087: imageROM = 8'd79;
                3088: imageROM = 8'd20;
                3089: imageROM = 8'd70;
                3090: imageROM = 8'd130;
                3091: imageROM = 8'd73;
                3092: imageROM = 8'd191;
                3093: imageROM = 8'd143;
                3094: imageROM = 8'd79;
                3095: imageROM = 8'd19;
                3096: imageROM = 8'd69;
                3097: imageROM = 8'd132;
                3098: imageROM = 8'd73;
                3099: imageROM = 8'd191;
                3100: imageROM = 8'd143;
                3101: imageROM = 8'd78;
                3102: imageROM = 8'd18;
                3103: imageROM = 8'd70;
                3104: imageROM = 8'd132;
                3105: imageROM = 8'd74;
                3106: imageROM = 8'd191;
                3107: imageROM = 8'd144;
                3108: imageROM = 8'd77;
                3109: imageROM = 8'd16;
                3110: imageROM = 8'd70;
                3111: imageROM = 8'd133;
                3112: imageROM = 8'd75;
                3113: imageROM = 8'd191;
                3114: imageROM = 8'd145;
                3115: imageROM = 8'd75;
                3116: imageROM = 8'd16;
                3117: imageROM = 8'd70;
                3118: imageROM = 8'd133;
                3119: imageROM = 8'd82;
                3120: imageROM = 8'd191;
                3121: imageROM = 8'd139;
                3122: imageROM = 8'd74;
                3123: imageROM = 8'd15;
                3124: imageROM = 8'd70;
                3125: imageROM = 8'd135;
                3126: imageROM = 8'd81;
                3127: imageROM = 8'd191;
                3128: imageROM = 8'd140;
                3129: imageROM = 8'd73;
                3130: imageROM = 8'd15;
                3131: imageROM = 8'd69;
                3132: imageROM = 8'd137;
                3133: imageROM = 8'd79;
                3134: imageROM = 8'd191;
                3135: imageROM = 8'd142;
                3136: imageROM = 8'd72;
                3137: imageROM = 8'd14;
                3138: imageROM = 8'd70;
                3139: imageROM = 8'd138;
                3140: imageROM = 8'd77;
                3141: imageROM = 8'd191;
                3142: imageROM = 8'd144;
                3143: imageROM = 8'd71;
                3144: imageROM = 8'd13;
                3145: imageROM = 8'd70;
                3146: imageROM = 8'd141;
                3147: imageROM = 8'd74;
                3148: imageROM = 8'd191;
                3149: imageROM = 8'd145;
                3150: imageROM = 8'd71;
                3151: imageROM = 8'd13;
                3152: imageROM = 8'd70;
                3153: imageROM = 8'd144;
                3154: imageROM = 8'd70;
                3155: imageROM = 8'd191;
                3156: imageROM = 8'd146;
                3157: imageROM = 8'd70;
                3158: imageROM = 8'd13;
                3159: imageROM = 8'd70;
                3160: imageROM = 8'd191;
                3161: imageROM = 8'd169;
                3162: imageROM = 8'd70;
                3163: imageROM = 8'd13;
                3164: imageROM = 8'd70;
                3165: imageROM = 8'd191;
                3166: imageROM = 8'd168;
                3167: imageROM = 8'd71;
                3168: imageROM = 8'd12;
                3169: imageROM = 8'd70;
                3170: imageROM = 8'd191;
                3171: imageROM = 8'd169;
                3172: imageROM = 8'd71;
                3173: imageROM = 8'd12;
                3174: imageROM = 8'd70;
                3175: imageROM = 8'd191;
                3176: imageROM = 8'd169;
                3177: imageROM = 8'd70;
            // r06.bmp
                3178: imageROM = 8'd63;
                3179: imageROM = 8'd63;
                3180: imageROM = 8'd63;
                3181: imageROM = 8'd63;
                3182: imageROM = 8'd63;
                3183: imageROM = 8'd63;
                3184: imageROM = 8'd63;
                3185: imageROM = 8'd63;
                3186: imageROM = 8'd63;
                3187: imageROM = 8'd63;
                3188: imageROM = 8'd63;
                3189: imageROM = 8'd63;
                3190: imageROM = 8'd63;
                3191: imageROM = 8'd63;
                3192: imageROM = 8'd63;
                3193: imageROM = 8'd63;
                3194: imageROM = 8'd63;
                3195: imageROM = 8'd63;
                3196: imageROM = 8'd63;
                3197: imageROM = 8'd63;
                3198: imageROM = 8'd63;
                3199: imageROM = 8'd63;
                3200: imageROM = 8'd63;
                3201: imageROM = 8'd63;
                3202: imageROM = 8'd63;
                3203: imageROM = 8'd63;
                3204: imageROM = 8'd63;
                3205: imageROM = 8'd63;
                3206: imageROM = 8'd62;
                3207: imageROM = 8'd79;
                3208: imageROM = 8'd63;
                3209: imageROM = 8'd46;
                3210: imageROM = 8'd88;
                3211: imageROM = 8'd63;
                3212: imageROM = 8'd38;
                3213: imageROM = 8'd94;
                3214: imageROM = 8'd63;
                3215: imageROM = 8'd34;
                3216: imageROM = 8'd97;
                3217: imageROM = 8'd63;
                3218: imageROM = 8'd30;
                3219: imageROM = 8'd101;
                3220: imageROM = 8'd63;
                3221: imageROM = 8'd26;
                3222: imageROM = 8'd104;
                3223: imageROM = 8'd63;
                3224: imageROM = 8'd24;
                3225: imageROM = 8'd75;
                3226: imageROM = 8'd147;
                3227: imageROM = 8'd77;
                3228: imageROM = 8'd63;
                3229: imageROM = 8'd20;
                3230: imageROM = 8'd74;
                3231: imageROM = 8'd154;
                3232: imageROM = 8'd74;
                3233: imageROM = 8'd63;
                3234: imageROM = 8'd18;
                3235: imageROM = 8'd73;
                3236: imageROM = 8'd158;
                3237: imageROM = 8'd73;
                3238: imageROM = 8'd63;
                3239: imageROM = 8'd16;
                3240: imageROM = 8'd73;
                3241: imageROM = 8'd161;
                3242: imageROM = 8'd72;
                3243: imageROM = 8'd63;
                3244: imageROM = 8'd14;
                3245: imageROM = 8'd72;
                3246: imageROM = 8'd164;
                3247: imageROM = 8'd72;
                3248: imageROM = 8'd63;
                3249: imageROM = 8'd12;
                3250: imageROM = 8'd72;
                3251: imageROM = 8'd166;
                3252: imageROM = 8'd71;
                3253: imageROM = 8'd63;
                3254: imageROM = 8'd11;
                3255: imageROM = 8'd72;
                3256: imageROM = 8'd168;
                3257: imageROM = 8'd71;
                3258: imageROM = 8'd63;
                3259: imageROM = 8'd9;
                3260: imageROM = 8'd72;
                3261: imageROM = 8'd170;
                3262: imageROM = 8'd71;
                3263: imageROM = 8'd63;
                3264: imageROM = 8'd7;
                3265: imageROM = 8'd72;
                3266: imageROM = 8'd135;
                3267: imageROM = 8'd67;
                3268: imageROM = 8'd162;
                3269: imageROM = 8'd70;
                3270: imageROM = 8'd63;
                3271: imageROM = 8'd6;
                3272: imageROM = 8'd72;
                3273: imageROM = 8'd134;
                3274: imageROM = 8'd71;
                3275: imageROM = 8'd160;
                3276: imageROM = 8'd71;
                3277: imageROM = 8'd63;
                3278: imageROM = 8'd5;
                3279: imageROM = 8'd71;
                3280: imageROM = 8'd134;
                3281: imageROM = 8'd72;
                3282: imageROM = 8'd159;
                3283: imageROM = 8'd72;
                3284: imageROM = 8'd63;
                3285: imageROM = 8'd4;
                3286: imageROM = 8'd71;
                3287: imageROM = 8'd135;
                3288: imageROM = 8'd73;
                3289: imageROM = 8'd145;
                3290: imageROM = 8'd69;
                3291: imageROM = 8'd135;
                3292: imageROM = 8'd74;
                3293: imageROM = 8'd63;
                3294: imageROM = 8'd2;
                3295: imageROM = 8'd71;
                3296: imageROM = 8'd136;
                3297: imageROM = 8'd74;
                3298: imageROM = 8'd141;
                3299: imageROM = 8'd75;
                3300: imageROM = 8'd132;
                3301: imageROM = 8'd74;
                3302: imageROM = 8'd63;
                3303: imageROM = 8'd1;
                3304: imageROM = 8'd71;
                3305: imageROM = 8'd137;
                3306: imageROM = 8'd74;
                3307: imageROM = 8'd139;
                3308: imageROM = 8'd78;
                3309: imageROM = 8'd131;
                3310: imageROM = 8'd75;
                3311: imageROM = 8'd63;
                3312: imageROM = 8'd70;
                3313: imageROM = 8'd138;
                3314: imageROM = 8'd74;
                3315: imageROM = 8'd138;
                3316: imageROM = 8'd80;
                3317: imageROM = 8'd130;
                3318: imageROM = 8'd75;
                3319: imageROM = 8'd62;
                3320: imageROM = 8'd71;
                3321: imageROM = 8'd138;
                3322: imageROM = 8'd74;
                3323: imageROM = 8'd137;
                3324: imageROM = 8'd82;
                3325: imageROM = 8'd129;
                3326: imageROM = 8'd75;
                3327: imageROM = 8'd61;
                3328: imageROM = 8'd71;
                3329: imageROM = 8'd139;
                3330: imageROM = 8'd74;
                3331: imageROM = 8'd137;
                3332: imageROM = 8'd95;
                3333: imageROM = 8'd60;
                3334: imageROM = 8'd70;
                3335: imageROM = 8'd140;
                3336: imageROM = 8'd74;
                3337: imageROM = 8'd136;
                3338: imageROM = 8'd71;
                3339: imageROM = 8'd198;
                3340: imageROM = 8'd83;
                3341: imageROM = 8'd59;
                3342: imageROM = 8'd70;
                3343: imageROM = 8'd141;
                3344: imageROM = 8'd74;
                3345: imageROM = 8'd136;
                3346: imageROM = 8'd70;
                3347: imageROM = 8'd200;
                3348: imageROM = 8'd83;
                3349: imageROM = 8'd57;
                3350: imageROM = 8'd71;
                3351: imageROM = 8'd142;
                3352: imageROM = 8'd72;
                3353: imageROM = 8'd136;
                3354: imageROM = 8'd70;
                3355: imageROM = 8'd202;
                3356: imageROM = 8'd70;
                3357: imageROM = 8'd130;
                3358: imageROM = 8'd67;
                3359: imageROM = 8'd129;
                3360: imageROM = 8'd71;
                3361: imageROM = 8'd56;
                3362: imageROM = 8'd70;
                3363: imageROM = 8'd144;
                3364: imageROM = 8'd71;
                3365: imageROM = 8'd136;
                3366: imageROM = 8'd70;
                3367: imageROM = 8'd202;
                3368: imageROM = 8'd71;
                3369: imageROM = 8'd134;
                3370: imageROM = 8'd71;
                3371: imageROM = 8'd54;
                3372: imageROM = 8'd70;
                3373: imageROM = 8'd147;
                3374: imageROM = 8'd65;
                3375: imageROM = 8'd129;
                3376: imageROM = 8'd65;
                3377: imageROM = 8'd138;
                3378: imageROM = 8'd69;
                3379: imageROM = 8'd204;
                3380: imageROM = 8'd70;
                3381: imageROM = 8'd134;
                3382: imageROM = 8'd72;
                3383: imageROM = 8'd53;
                3384: imageROM = 8'd70;
                3385: imageROM = 8'd159;
                3386: imageROM = 8'd70;
                3387: imageROM = 8'd204;
                3388: imageROM = 8'd70;
                3389: imageROM = 8'd135;
                3390: imageROM = 8'd72;
                3391: imageROM = 8'd51;
                3392: imageROM = 8'd70;
                3393: imageROM = 8'd160;
                3394: imageROM = 8'd70;
                3395: imageROM = 8'd204;
                3396: imageROM = 8'd70;
                3397: imageROM = 8'd136;
                3398: imageROM = 8'd73;
                3399: imageROM = 8'd49;
                3400: imageROM = 8'd70;
                3401: imageROM = 8'd160;
                3402: imageROM = 8'd70;
                3403: imageROM = 8'd205;
                3404: imageROM = 8'd70;
                3405: imageROM = 8'd136;
                3406: imageROM = 8'd73;
                3407: imageROM = 8'd47;
                3408: imageROM = 8'd70;
                3409: imageROM = 8'd161;
                3410: imageROM = 8'd70;
                3411: imageROM = 8'd205;
                3412: imageROM = 8'd70;
                3413: imageROM = 8'd138;
                3414: imageROM = 8'd72;
                3415: imageROM = 8'd46;
                3416: imageROM = 8'd70;
                3417: imageROM = 8'd161;
                3418: imageROM = 8'd70;
                3419: imageROM = 8'd205;
                3420: imageROM = 8'd70;
                3421: imageROM = 8'd139;
                3422: imageROM = 8'd72;
                3423: imageROM = 8'd44;
                3424: imageROM = 8'd70;
                3425: imageROM = 8'd162;
                3426: imageROM = 8'd70;
                3427: imageROM = 8'd205;
                3428: imageROM = 8'd70;
                3429: imageROM = 8'd140;
                3430: imageROM = 8'd71;
                3431: imageROM = 8'd44;
                3432: imageROM = 8'd70;
                3433: imageROM = 8'd162;
                3434: imageROM = 8'd70;
                3435: imageROM = 8'd205;
                3436: imageROM = 8'd70;
                3437: imageROM = 8'd141;
                3438: imageROM = 8'd71;
                3439: imageROM = 8'd43;
                3440: imageROM = 8'd70;
                3441: imageROM = 8'd162;
                3442: imageROM = 8'd70;
                3443: imageROM = 8'd205;
                3444: imageROM = 8'd70;
                3445: imageROM = 8'd142;
                3446: imageROM = 8'd71;
                3447: imageROM = 8'd42;
                3448: imageROM = 8'd69;
                3449: imageROM = 8'd163;
                3450: imageROM = 8'd70;
                3451: imageROM = 8'd205;
                3452: imageROM = 8'd70;
                3453: imageROM = 8'd143;
                3454: imageROM = 8'd70;
                3455: imageROM = 8'd42;
                3456: imageROM = 8'd69;
                3457: imageROM = 8'd163;
                3458: imageROM = 8'd70;
                3459: imageROM = 8'd205;
                3460: imageROM = 8'd70;
                3461: imageROM = 8'd144;
                3462: imageROM = 8'd70;
                3463: imageROM = 8'd41;
                3464: imageROM = 8'd69;
                3465: imageROM = 8'd163;
                3466: imageROM = 8'd70;
                3467: imageROM = 8'd205;
                3468: imageROM = 8'd70;
                3469: imageROM = 8'd144;
                3470: imageROM = 8'd70;
                3471: imageROM = 8'd41;
                3472: imageROM = 8'd69;
                3473: imageROM = 8'd163;
                3474: imageROM = 8'd70;
                3475: imageROM = 8'd205;
                3476: imageROM = 8'd70;
                3477: imageROM = 8'd144;
                3478: imageROM = 8'd70;
                3479: imageROM = 8'd41;
                3480: imageROM = 8'd69;
                3481: imageROM = 8'd163;
                3482: imageROM = 8'd70;
                3483: imageROM = 8'd205;
                3484: imageROM = 8'd70;
                3485: imageROM = 8'd145;
                3486: imageROM = 8'd69;
                3487: imageROM = 8'd41;
                3488: imageROM = 8'd69;
                3489: imageROM = 8'd164;
                3490: imageROM = 8'd69;
                3491: imageROM = 8'd205;
                3492: imageROM = 8'd70;
                3493: imageROM = 8'd145;
                3494: imageROM = 8'd69;
                3495: imageROM = 8'd41;
                3496: imageROM = 8'd70;
                3497: imageROM = 8'd163;
                3498: imageROM = 8'd70;
                3499: imageROM = 8'd204;
                3500: imageROM = 8'd70;
                3501: imageROM = 8'd145;
                3502: imageROM = 8'd69;
                3503: imageROM = 8'd41;
                3504: imageROM = 8'd70;
                3505: imageROM = 8'd163;
                3506: imageROM = 8'd70;
                3507: imageROM = 8'd204;
                3508: imageROM = 8'd70;
                3509: imageROM = 8'd145;
                3510: imageROM = 8'd69;
                3511: imageROM = 8'd41;
                3512: imageROM = 8'd70;
                3513: imageROM = 8'd163;
                3514: imageROM = 8'd70;
                3515: imageROM = 8'd203;
                3516: imageROM = 8'd70;
                3517: imageROM = 8'd146;
                3518: imageROM = 8'd69;
                3519: imageROM = 8'd42;
                3520: imageROM = 8'd69;
                3521: imageROM = 8'd164;
                3522: imageROM = 8'd70;
                3523: imageROM = 8'd202;
                3524: imageROM = 8'd70;
                3525: imageROM = 8'd146;
                3526: imageROM = 8'd69;
                3527: imageROM = 8'd42;
                3528: imageROM = 8'd69;
                3529: imageROM = 8'd164;
                3530: imageROM = 8'd70;
                3531: imageROM = 8'd202;
                3532: imageROM = 8'd70;
                3533: imageROM = 8'd146;
                3534: imageROM = 8'd69;
                3535: imageROM = 8'd42;
                3536: imageROM = 8'd70;
                3537: imageROM = 8'd163;
                3538: imageROM = 8'd70;
                3539: imageROM = 8'd201;
                3540: imageROM = 8'd71;
                3541: imageROM = 8'd146;
                3542: imageROM = 8'd69;
                3543: imageROM = 8'd42;
                3544: imageROM = 8'd70;
                3545: imageROM = 8'd164;
                3546: imageROM = 8'd70;
                3547: imageROM = 8'd200;
                3548: imageROM = 8'd70;
                3549: imageROM = 8'd147;
                3550: imageROM = 8'd69;
                3551: imageROM = 8'd42;
                3552: imageROM = 8'd70;
                3553: imageROM = 8'd164;
                3554: imageROM = 8'd70;
                3555: imageROM = 8'd199;
                3556: imageROM = 8'd71;
                3557: imageROM = 8'd147;
                3558: imageROM = 8'd69;
                3559: imageROM = 8'd43;
                3560: imageROM = 8'd69;
                3561: imageROM = 8'd164;
                3562: imageROM = 8'd71;
                3563: imageROM = 8'd197;
                3564: imageROM = 8'd71;
                3565: imageROM = 8'd147;
                3566: imageROM = 8'd70;
                3567: imageROM = 8'd43;
                3568: imageROM = 8'd70;
                3569: imageROM = 8'd164;
                3570: imageROM = 8'd71;
                3571: imageROM = 8'd196;
                3572: imageROM = 8'd71;
                3573: imageROM = 8'd147;
                3574: imageROM = 8'd70;
                3575: imageROM = 8'd43;
                3576: imageROM = 8'd69;
                3577: imageROM = 8'd165;
                3578: imageROM = 8'd71;
                3579: imageROM = 8'd195;
                3580: imageROM = 8'd71;
                3581: imageROM = 8'd148;
                3582: imageROM = 8'd70;
                3583: imageROM = 8'd43;
                3584: imageROM = 8'd70;
                3585: imageROM = 8'd165;
                3586: imageROM = 8'd71;
                3587: imageROM = 8'd194;
                3588: imageROM = 8'd70;
                3589: imageROM = 8'd149;
                3590: imageROM = 8'd70;
                3591: imageROM = 8'd43;
                3592: imageROM = 8'd70;
                3593: imageROM = 8'd166;
                3594: imageROM = 8'd78;
                3595: imageROM = 8'd149;
                3596: imageROM = 8'd70;
                3597: imageROM = 8'd43;
                3598: imageROM = 8'd70;
                3599: imageROM = 8'd167;
                3600: imageROM = 8'd76;
                3601: imageROM = 8'd150;
                3602: imageROM = 8'd70;
                3603: imageROM = 8'd43;
                3604: imageROM = 8'd70;
                3605: imageROM = 8'd167;
                3606: imageROM = 8'd75;
                3607: imageROM = 8'd151;
                3608: imageROM = 8'd70;
                3609: imageROM = 8'd43;
                3610: imageROM = 8'd70;
                3611: imageROM = 8'd168;
                3612: imageROM = 8'd74;
                3613: imageROM = 8'd151;
                3614: imageROM = 8'd70;
                3615: imageROM = 8'd43;
                3616: imageROM = 8'd70;
                3617: imageROM = 8'd169;
                3618: imageROM = 8'd72;
                3619: imageROM = 8'd152;
                3620: imageROM = 8'd70;
                3621: imageROM = 8'd43;
                3622: imageROM = 8'd71;
                3623: imageROM = 8'd168;
                3624: imageROM = 8'd72;
                3625: imageROM = 8'd152;
                3626: imageROM = 8'd70;
                3627: imageROM = 8'd43;
                3628: imageROM = 8'd71;
                3629: imageROM = 8'd169;
                3630: imageROM = 8'd70;
                3631: imageROM = 8'd153;
                3632: imageROM = 8'd70;
                3633: imageROM = 8'd43;
                3634: imageROM = 8'd71;
                3635: imageROM = 8'd170;
                3636: imageROM = 8'd69;
                3637: imageROM = 8'd153;
                3638: imageROM = 8'd70;
                3639: imageROM = 8'd43;
                3640: imageROM = 8'd72;
                3641: imageROM = 8'd170;
                3642: imageROM = 8'd67;
                3643: imageROM = 8'd155;
                3644: imageROM = 8'd69;
                3645: imageROM = 8'd43;
                3646: imageROM = 8'd72;
                3647: imageROM = 8'd170;
                3648: imageROM = 8'd67;
                3649: imageROM = 8'd155;
                3650: imageROM = 8'd70;
                3651: imageROM = 8'd41;
                3652: imageROM = 8'd74;
                3653: imageROM = 8'd170;
                3654: imageROM = 8'd65;
                3655: imageROM = 8'd156;
                3656: imageROM = 8'd71;
                3657: imageROM = 8'd40;
                3658: imageROM = 8'd74;
                3659: imageROM = 8'd191;
                3660: imageROM = 8'd137;
                3661: imageROM = 8'd71;
                3662: imageROM = 8'd39;
                3663: imageROM = 8'd75;
                3664: imageROM = 8'd191;
                3665: imageROM = 8'd136;
                3666: imageROM = 8'd72;
                3667: imageROM = 8'd38;
                3668: imageROM = 8'd75;
                3669: imageROM = 8'd191;
                3670: imageROM = 8'd137;
                3671: imageROM = 8'd72;
                3672: imageROM = 8'd37;
                3673: imageROM = 8'd76;
                3674: imageROM = 8'd191;
                3675: imageROM = 8'd137;
                3676: imageROM = 8'd72;
                3677: imageROM = 8'd36;
                3678: imageROM = 8'd69;
                3679: imageROM = 8'd1;
                3680: imageROM = 8'd71;
                3681: imageROM = 8'd191;
                3682: imageROM = 8'd137;
                3683: imageROM = 8'd72;
                3684: imageROM = 8'd35;
                3685: imageROM = 8'd70;
                3686: imageROM = 8'd129;
                3687: imageROM = 8'd71;
                3688: imageROM = 8'd191;
                3689: imageROM = 8'd137;
                3690: imageROM = 8'd72;
                3691: imageROM = 8'd34;
                3692: imageROM = 8'd70;
                3693: imageROM = 8'd130;
                3694: imageROM = 8'd70;
                3695: imageROM = 8'd191;
                3696: imageROM = 8'd138;
                3697: imageROM = 8'd73;
                3698: imageROM = 8'd32;
                3699: imageROM = 8'd69;
                3700: imageROM = 8'd132;
                3701: imageROM = 8'd70;
                3702: imageROM = 8'd191;
                3703: imageROM = 8'd138;
                3704: imageROM = 8'd73;
                3705: imageROM = 8'd31;
                3706: imageROM = 8'd69;
                3707: imageROM = 8'd133;
                3708: imageROM = 8'd70;
                3709: imageROM = 8'd191;
                3710: imageROM = 8'd138;
                3711: imageROM = 8'd73;
                3712: imageROM = 8'd30;
                3713: imageROM = 8'd69;
                3714: imageROM = 8'd133;
                3715: imageROM = 8'd71;
                3716: imageROM = 8'd191;
                3717: imageROM = 8'd139;
                3718: imageROM = 8'd73;
                3719: imageROM = 8'd28;
                3720: imageROM = 8'd69;
                3721: imageROM = 8'd134;
                3722: imageROM = 8'd71;
                3723: imageROM = 8'd191;
                3724: imageROM = 8'd139;
                3725: imageROM = 8'd73;
                3726: imageROM = 8'd27;
                3727: imageROM = 8'd69;
                3728: imageROM = 8'd135;
                3729: imageROM = 8'd72;
                3730: imageROM = 8'd191;
                3731: imageROM = 8'd138;
                3732: imageROM = 8'd74;
                3733: imageROM = 8'd25;
                3734: imageROM = 8'd69;
                3735: imageROM = 8'd136;
                3736: imageROM = 8'd72;
                3737: imageROM = 8'd191;
                3738: imageROM = 8'd138;
                3739: imageROM = 8'd74;
                3740: imageROM = 8'd24;
                3741: imageROM = 8'd69;
                3742: imageROM = 8'd137;
                3743: imageROM = 8'd73;
                3744: imageROM = 8'd191;
                3745: imageROM = 8'd138;
                3746: imageROM = 8'd74;
                3747: imageROM = 8'd22;
                3748: imageROM = 8'd69;
                3749: imageROM = 8'd138;
                3750: imageROM = 8'd73;
                3751: imageROM = 8'd191;
                3752: imageROM = 8'd138;
                3753: imageROM = 8'd75;
                3754: imageROM = 8'd20;
                3755: imageROM = 8'd70;
                3756: imageROM = 8'd139;
                3757: imageROM = 8'd73;
                3758: imageROM = 8'd191;
                3759: imageROM = 8'd138;
                3760: imageROM = 8'd74;
                3761: imageROM = 8'd19;
                3762: imageROM = 8'd70;
                3763: imageROM = 8'd140;
                3764: imageROM = 8'd75;
                3765: imageROM = 8'd191;
                3766: imageROM = 8'd137;
                3767: imageROM = 8'd74;
                3768: imageROM = 8'd17;
                3769: imageROM = 8'd70;
                3770: imageROM = 8'd141;
                3771: imageROM = 8'd82;
                3772: imageROM = 8'd191;
                3773: imageROM = 8'd130;
                3774: imageROM = 8'd75;
                3775: imageROM = 8'd16;
                3776: imageROM = 8'd70;
                3777: imageROM = 8'd142;
                3778: imageROM = 8'd81;
                3779: imageROM = 8'd191;
                3780: imageROM = 8'd131;
                3781: imageROM = 8'd74;
                3782: imageROM = 8'd15;
                3783: imageROM = 8'd70;
                3784: imageROM = 8'd144;
                3785: imageROM = 8'd79;
                3786: imageROM = 8'd191;
                3787: imageROM = 8'd133;
                3788: imageROM = 8'd73;
            // r07.bmp
                3789: imageROM = 8'd63;
                3790: imageROM = 8'd63;
                3791: imageROM = 8'd63;
                3792: imageROM = 8'd63;
                3793: imageROM = 8'd63;
                3794: imageROM = 8'd63;
                3795: imageROM = 8'd63;
                3796: imageROM = 8'd63;
                3797: imageROM = 8'd63;
                3798: imageROM = 8'd63;
                3799: imageROM = 8'd63;
                3800: imageROM = 8'd63;
                3801: imageROM = 8'd63;
                3802: imageROM = 8'd63;
                3803: imageROM = 8'd63;
                3804: imageROM = 8'd63;
                3805: imageROM = 8'd63;
                3806: imageROM = 8'd63;
                3807: imageROM = 8'd63;
                3808: imageROM = 8'd63;
                3809: imageROM = 8'd63;
                3810: imageROM = 8'd63;
                3811: imageROM = 8'd63;
                3812: imageROM = 8'd63;
                3813: imageROM = 8'd63;
                3814: imageROM = 8'd63;
                3815: imageROM = 8'd63;
                3816: imageROM = 8'd63;
                3817: imageROM = 8'd63;
                3818: imageROM = 8'd63;
                3819: imageROM = 8'd63;
                3820: imageROM = 8'd63;
                3821: imageROM = 8'd63;
                3822: imageROM = 8'd63;
                3823: imageROM = 8'd63;
                3824: imageROM = 8'd63;
                3825: imageROM = 8'd63;
                3826: imageROM = 8'd63;
                3827: imageROM = 8'd63;
                3828: imageROM = 8'd63;
                3829: imageROM = 8'd63;
                3830: imageROM = 8'd22;
                3831: imageROM = 8'd85;
                3832: imageROM = 8'd63;
                3833: imageROM = 8'd40;
                3834: imageROM = 8'd93;
                3835: imageROM = 8'd63;
                3836: imageROM = 8'd33;
                3837: imageROM = 8'd98;
                3838: imageROM = 8'd63;
                3839: imageROM = 8'd29;
                3840: imageROM = 8'd102;
                3841: imageROM = 8'd63;
                3842: imageROM = 8'd25;
                3843: imageROM = 8'd105;
                3844: imageROM = 8'd63;
                3845: imageROM = 8'd23;
                3846: imageROM = 8'd78;
                3847: imageROM = 8'd144;
                3848: imageROM = 8'd77;
                3849: imageROM = 8'd63;
                3850: imageROM = 8'd20;
                3851: imageROM = 8'd76;
                3852: imageROM = 8'd152;
                3853: imageROM = 8'd74;
                3854: imageROM = 8'd63;
                3855: imageROM = 8'd18;
                3856: imageROM = 8'd74;
                3857: imageROM = 8'd158;
                3858: imageROM = 8'd72;
                3859: imageROM = 8'd63;
                3860: imageROM = 8'd15;
                3861: imageROM = 8'd74;
                3862: imageROM = 8'd162;
                3863: imageROM = 8'd71;
                3864: imageROM = 8'd63;
                3865: imageROM = 8'd13;
                3866: imageROM = 8'd73;
                3867: imageROM = 8'd165;
                3868: imageROM = 8'd71;
                3869: imageROM = 8'd63;
                3870: imageROM = 8'd11;
                3871: imageROM = 8'd73;
                3872: imageROM = 8'd167;
                3873: imageROM = 8'd71;
                3874: imageROM = 8'd63;
                3875: imageROM = 8'd9;
                3876: imageROM = 8'd72;
                3877: imageROM = 8'd170;
                3878: imageROM = 8'd70;
                3879: imageROM = 8'd63;
                3880: imageROM = 8'd8;
                3881: imageROM = 8'd72;
                3882: imageROM = 8'd172;
                3883: imageROM = 8'd70;
                3884: imageROM = 8'd63;
                3885: imageROM = 8'd6;
                3886: imageROM = 8'd72;
                3887: imageROM = 8'd173;
                3888: imageROM = 8'd71;
                3889: imageROM = 8'd63;
                3890: imageROM = 8'd4;
                3891: imageROM = 8'd71;
                3892: imageROM = 8'd176;
                3893: imageROM = 8'd70;
                3894: imageROM = 8'd63;
                3895: imageROM = 8'd3;
                3896: imageROM = 8'd71;
                3897: imageROM = 8'd178;
                3898: imageROM = 8'd70;
                3899: imageROM = 8'd63;
                3900: imageROM = 8'd1;
                3901: imageROM = 8'd71;
                3902: imageROM = 8'd141;
                3903: imageROM = 8'd68;
                3904: imageROM = 8'd162;
                3905: imageROM = 8'd70;
                3906: imageROM = 8'd63;
                3907: imageROM = 8'd71;
                3908: imageROM = 8'd140;
                3909: imageROM = 8'd72;
                3910: imageROM = 8'd159;
                3911: imageROM = 8'd72;
                3912: imageROM = 8'd61;
                3913: imageROM = 8'd71;
                3914: imageROM = 8'd141;
                3915: imageROM = 8'd72;
                3916: imageROM = 8'd158;
                3917: imageROM = 8'd73;
                3918: imageROM = 8'd60;
                3919: imageROM = 8'd71;
                3920: imageROM = 8'd142;
                3921: imageROM = 8'd73;
                3922: imageROM = 8'd157;
                3923: imageROM = 8'd74;
                3924: imageROM = 8'd58;
                3925: imageROM = 8'd71;
                3926: imageROM = 8'd142;
                3927: imageROM = 8'd74;
                3928: imageROM = 8'd141;
                3929: imageROM = 8'd72;
                3930: imageROM = 8'd135;
                3931: imageROM = 8'd75;
                3932: imageROM = 8'd57;
                3933: imageROM = 8'd71;
                3934: imageROM = 8'd143;
                3935: imageROM = 8'd75;
                3936: imageROM = 8'd138;
                3937: imageROM = 8'd76;
                3938: imageROM = 8'd133;
                3939: imageROM = 8'd76;
                3940: imageROM = 8'd56;
                3941: imageROM = 8'd70;
                3942: imageROM = 8'd144;
                3943: imageROM = 8'd75;
                3944: imageROM = 8'd137;
                3945: imageROM = 8'd78;
                3946: imageROM = 8'd132;
                3947: imageROM = 8'd77;
                3948: imageROM = 8'd54;
                3949: imageROM = 8'd71;
                3950: imageROM = 8'd144;
                3951: imageROM = 8'd75;
                3952: imageROM = 8'd136;
                3953: imageROM = 8'd80;
                3954: imageROM = 8'd131;
                3955: imageROM = 8'd77;
                3956: imageROM = 8'd53;
                3957: imageROM = 8'd71;
                3958: imageROM = 8'd145;
                3959: imageROM = 8'd75;
                3960: imageROM = 8'd135;
                3961: imageROM = 8'd82;
                3962: imageROM = 8'd131;
                3963: imageROM = 8'd77;
                3964: imageROM = 8'd52;
                3965: imageROM = 8'd70;
                3966: imageROM = 8'd147;
                3967: imageROM = 8'd74;
                3968: imageROM = 8'd135;
                3969: imageROM = 8'd83;
                3970: imageROM = 8'd131;
                3971: imageROM = 8'd77;
                3972: imageROM = 8'd50;
                3973: imageROM = 8'd70;
                3974: imageROM = 8'd148;
                3975: imageROM = 8'd73;
                3976: imageROM = 8'd135;
                3977: imageROM = 8'd71;
                3978: imageROM = 8'd199;
                3979: imageROM = 8'd70;
                3980: imageROM = 8'd131;
                3981: imageROM = 8'd70;
                3982: imageROM = 8'd129;
                3983: imageROM = 8'd70;
                3984: imageROM = 8'd50;
                3985: imageROM = 8'd70;
                3986: imageROM = 8'd149;
                3987: imageROM = 8'd72;
                3988: imageROM = 8'd135;
                3989: imageROM = 8'd70;
                3990: imageROM = 8'd200;
                3991: imageROM = 8'd71;
                3992: imageROM = 8'd132;
                3993: imageROM = 8'd66;
                3994: imageROM = 8'd131;
                3995: imageROM = 8'd71;
                3996: imageROM = 8'd48;
                3997: imageROM = 8'd70;
                3998: imageROM = 8'd151;
                3999: imageROM = 8'd70;
                4000: imageROM = 8'd135;
                4001: imageROM = 8'd70;
                4002: imageROM = 8'd202;
                4003: imageROM = 8'd70;
                4004: imageROM = 8'd138;
                4005: imageROM = 8'd71;
                4006: imageROM = 8'd47;
                4007: imageROM = 8'd70;
                4008: imageROM = 8'd164;
                4009: imageROM = 8'd70;
                4010: imageROM = 8'd203;
                4011: imageROM = 8'd70;
                4012: imageROM = 8'd138;
                4013: imageROM = 8'd70;
                4014: imageROM = 8'd46;
                4015: imageROM = 8'd70;
                4016: imageROM = 8'd165;
                4017: imageROM = 8'd69;
                4018: imageROM = 8'd204;
                4019: imageROM = 8'd70;
                4020: imageROM = 8'd139;
                4021: imageROM = 8'd70;
                4022: imageROM = 8'd45;
                4023: imageROM = 8'd70;
                4024: imageROM = 8'd164;
                4025: imageROM = 8'd70;
                4026: imageROM = 8'd204;
                4027: imageROM = 8'd70;
                4028: imageROM = 8'd139;
                4029: imageROM = 8'd70;
                4030: imageROM = 8'd44;
                4031: imageROM = 8'd70;
                4032: imageROM = 8'd165;
                4033: imageROM = 8'd70;
                4034: imageROM = 8'd205;
                4035: imageROM = 8'd69;
                4036: imageROM = 8'd140;
                4037: imageROM = 8'd70;
                4038: imageROM = 8'd43;
                4039: imageROM = 8'd70;
                4040: imageROM = 8'd165;
                4041: imageROM = 8'd70;
                4042: imageROM = 8'd205;
                4043: imageROM = 8'd70;
                4044: imageROM = 8'd139;
                4045: imageROM = 8'd70;
                4046: imageROM = 8'd43;
                4047: imageROM = 8'd70;
                4048: imageROM = 8'd165;
                4049: imageROM = 8'd70;
                4050: imageROM = 8'd205;
                4051: imageROM = 8'd70;
                4052: imageROM = 8'd140;
                4053: imageROM = 8'd70;
                4054: imageROM = 8'd42;
                4055: imageROM = 8'd69;
                4056: imageROM = 8'd166;
                4057: imageROM = 8'd70;
                4058: imageROM = 8'd205;
                4059: imageROM = 8'd70;
                4060: imageROM = 8'd140;
                4061: imageROM = 8'd70;
                4062: imageROM = 8'd41;
                4063: imageROM = 8'd70;
                4064: imageROM = 8'd166;
                4065: imageROM = 8'd70;
                4066: imageROM = 8'd205;
                4067: imageROM = 8'd70;
                4068: imageROM = 8'd141;
                4069: imageROM = 8'd69;
                4070: imageROM = 8'd41;
                4071: imageROM = 8'd70;
                4072: imageROM = 8'd166;
                4073: imageROM = 8'd70;
                4074: imageROM = 8'd205;
                4075: imageROM = 8'd70;
                4076: imageROM = 8'd141;
                4077: imageROM = 8'd70;
                4078: imageROM = 8'd40;
                4079: imageROM = 8'd70;
                4080: imageROM = 8'd166;
                4081: imageROM = 8'd70;
                4082: imageROM = 8'd205;
                4083: imageROM = 8'd70;
                4084: imageROM = 8'd141;
                4085: imageROM = 8'd70;
                4086: imageROM = 8'd40;
                4087: imageROM = 8'd70;
                4088: imageROM = 8'd166;
                4089: imageROM = 8'd70;
                4090: imageROM = 8'd205;
                4091: imageROM = 8'd70;
                4092: imageROM = 8'd142;
                4093: imageROM = 8'd69;
                4094: imageROM = 8'd40;
                4095: imageROM = 8'd70;
                4096: imageROM = 8'd166;
                4097: imageROM = 8'd70;
                4098: imageROM = 8'd205;
                4099: imageROM = 8'd70;
                4100: imageROM = 8'd142;
                4101: imageROM = 8'd69;
                4102: imageROM = 8'd40;
                4103: imageROM = 8'd69;
                4104: imageROM = 8'd167;
                4105: imageROM = 8'd70;
                4106: imageROM = 8'd205;
                4107: imageROM = 8'd70;
                4108: imageROM = 8'd142;
                4109: imageROM = 8'd70;
                4110: imageROM = 8'd39;
                4111: imageROM = 8'd70;
                4112: imageROM = 8'd166;
                4113: imageROM = 8'd70;
                4114: imageROM = 8'd205;
                4115: imageROM = 8'd70;
                4116: imageROM = 8'd142;
                4117: imageROM = 8'd70;
                4118: imageROM = 8'd39;
                4119: imageROM = 8'd70;
                4120: imageROM = 8'd166;
                4121: imageROM = 8'd70;
                4122: imageROM = 8'd205;
                4123: imageROM = 8'd70;
                4124: imageROM = 8'd142;
                4125: imageROM = 8'd70;
                4126: imageROM = 8'd39;
                4127: imageROM = 8'd70;
                4128: imageROM = 8'd167;
                4129: imageROM = 8'd69;
                4130: imageROM = 8'd205;
                4131: imageROM = 8'd70;
                4132: imageROM = 8'd143;
                4133: imageROM = 8'd69;
                4134: imageROM = 8'd39;
                4135: imageROM = 8'd70;
                4136: imageROM = 8'd167;
                4137: imageROM = 8'd70;
                4138: imageROM = 8'd204;
                4139: imageROM = 8'd70;
                4140: imageROM = 8'd143;
                4141: imageROM = 8'd69;
                4142: imageROM = 8'd39;
                4143: imageROM = 8'd70;
                4144: imageROM = 8'd167;
                4145: imageROM = 8'd70;
                4146: imageROM = 8'd204;
                4147: imageROM = 8'd70;
                4148: imageROM = 8'd143;
                4149: imageROM = 8'd70;
                4150: imageROM = 8'd38;
                4151: imageROM = 8'd70;
                4152: imageROM = 8'd167;
                4153: imageROM = 8'd70;
                4154: imageROM = 8'd204;
                4155: imageROM = 8'd69;
                4156: imageROM = 8'd144;
                4157: imageROM = 8'd70;
                4158: imageROM = 8'd38;
                4159: imageROM = 8'd70;
                4160: imageROM = 8'd168;
                4161: imageROM = 8'd69;
                4162: imageROM = 8'd203;
                4163: imageROM = 8'd70;
                4164: imageROM = 8'd144;
                4165: imageROM = 8'd70;
                4166: imageROM = 8'd38;
                4167: imageROM = 8'd70;
                4168: imageROM = 8'd168;
                4169: imageROM = 8'd70;
                4170: imageROM = 8'd202;
                4171: imageROM = 8'd70;
                4172: imageROM = 8'd144;
                4173: imageROM = 8'd70;
                4174: imageROM = 8'd38;
                4175: imageROM = 8'd71;
                4176: imageROM = 8'd167;
                4177: imageROM = 8'd70;
                4178: imageROM = 8'd202;
                4179: imageROM = 8'd70;
                4180: imageROM = 8'd144;
                4181: imageROM = 8'd70;
                4182: imageROM = 8'd38;
                4183: imageROM = 8'd71;
                4184: imageROM = 8'd168;
                4185: imageROM = 8'd70;
                4186: imageROM = 8'd200;
                4187: imageROM = 8'd70;
                4188: imageROM = 8'd145;
                4189: imageROM = 8'd70;
                4190: imageROM = 8'd38;
                4191: imageROM = 8'd71;
                4192: imageROM = 8'd168;
                4193: imageROM = 8'd70;
                4194: imageROM = 8'd199;
                4195: imageROM = 8'd71;
                4196: imageROM = 8'd145;
                4197: imageROM = 8'd70;
                4198: imageROM = 8'd38;
                4199: imageROM = 8'd71;
                4200: imageROM = 8'd168;
                4201: imageROM = 8'd71;
                4202: imageROM = 8'd197;
                4203: imageROM = 8'd71;
                4204: imageROM = 8'd146;
                4205: imageROM = 8'd70;
                4206: imageROM = 8'd38;
                4207: imageROM = 8'd72;
                4208: imageROM = 8'd168;
                4209: imageROM = 8'd71;
                4210: imageROM = 8'd196;
                4211: imageROM = 8'd70;
                4212: imageROM = 8'd147;
                4213: imageROM = 8'd70;
                4214: imageROM = 8'd38;
                4215: imageROM = 8'd72;
                4216: imageROM = 8'd169;
                4217: imageROM = 8'd70;
                4218: imageROM = 8'd195;
                4219: imageROM = 8'd71;
                4220: imageROM = 8'd147;
                4221: imageROM = 8'd70;
                4222: imageROM = 8'd38;
                4223: imageROM = 8'd73;
                4224: imageROM = 8'd168;
                4225: imageROM = 8'd71;
                4226: imageROM = 8'd194;
                4227: imageROM = 8'd70;
                4228: imageROM = 8'd148;
                4229: imageROM = 8'd70;
                4230: imageROM = 8'd38;
                4231: imageROM = 8'd73;
                4232: imageROM = 8'd169;
                4233: imageROM = 8'd78;
                4234: imageROM = 8'd147;
                4235: imageROM = 8'd70;
                4236: imageROM = 8'd38;
                4237: imageROM = 8'd75;
                4238: imageROM = 8'd169;
                4239: imageROM = 8'd76;
                4240: imageROM = 8'd148;
                4241: imageROM = 8'd70;
                4242: imageROM = 8'd38;
                4243: imageROM = 8'd75;
                4244: imageROM = 8'd170;
                4245: imageROM = 8'd75;
                4246: imageROM = 8'd147;
                4247: imageROM = 8'd70;
                4248: imageROM = 8'd39;
                4249: imageROM = 8'd76;
                4250: imageROM = 8'd169;
                4251: imageROM = 8'd74;
                4252: imageROM = 8'd147;
                4253: imageROM = 8'd71;
                4254: imageROM = 8'd39;
                4255: imageROM = 8'd69;
                4256: imageROM = 8'd129;
                4257: imageROM = 8'd70;
                4258: imageROM = 8'd170;
                4259: imageROM = 8'd72;
                4260: imageROM = 8'd148;
                4261: imageROM = 8'd70;
                4262: imageROM = 8'd39;
                4263: imageROM = 8'd70;
                4264: imageROM = 8'd130;
                4265: imageROM = 8'd70;
                4266: imageROM = 8'd170;
                4267: imageROM = 8'd71;
                4268: imageROM = 8'd147;
                4269: imageROM = 8'd70;
                4270: imageROM = 8'd40;
                4271: imageROM = 8'd70;
                4272: imageROM = 8'd131;
                4273: imageROM = 8'd70;
                4274: imageROM = 8'd169;
                4275: imageROM = 8'd70;
                4276: imageROM = 8'd147;
                4277: imageROM = 8'd71;
                4278: imageROM = 8'd40;
                4279: imageROM = 8'd69;
                4280: imageROM = 8'd132;
                4281: imageROM = 8'd71;
                4282: imageROM = 8'd169;
                4283: imageROM = 8'd69;
                4284: imageROM = 8'd146;
                4285: imageROM = 8'd71;
                4286: imageROM = 8'd40;
                4287: imageROM = 8'd70;
                4288: imageROM = 8'd133;
                4289: imageROM = 8'd70;
                4290: imageROM = 8'd170;
                4291: imageROM = 8'd67;
                4292: imageROM = 8'd147;
                4293: imageROM = 8'd70;
                4294: imageROM = 8'd41;
                4295: imageROM = 8'd70;
                4296: imageROM = 8'd134;
                4297: imageROM = 8'd70;
                4298: imageROM = 8'd170;
                4299: imageROM = 8'd66;
                4300: imageROM = 8'd146;
                4301: imageROM = 8'd71;
                4302: imageROM = 8'd40;
                4303: imageROM = 8'd70;
                4304: imageROM = 8'd136;
                4305: imageROM = 8'd70;
                4306: imageROM = 8'd169;
                4307: imageROM = 8'd65;
                4308: imageROM = 8'd147;
                4309: imageROM = 8'd70;
                4310: imageROM = 8'd41;
                4311: imageROM = 8'd70;
                4312: imageROM = 8'd136;
                4313: imageROM = 8'd71;
                4314: imageROM = 8'd188;
                4315: imageROM = 8'd69;
                4316: imageROM = 8'd41;
                4317: imageROM = 8'd70;
                4318: imageROM = 8'd138;
                4319: imageROM = 8'd72;
                4320: imageROM = 8'd186;
                4321: imageROM = 8'd69;
                4322: imageROM = 8'd41;
                4323: imageROM = 8'd70;
                4324: imageROM = 8'd139;
                4325: imageROM = 8'd72;
                4326: imageROM = 8'd185;
                4327: imageROM = 8'd69;
                4328: imageROM = 8'd40;
                4329: imageROM = 8'd70;
                4330: imageROM = 8'd141;
                4331: imageROM = 8'd72;
                4332: imageROM = 8'd184;
                4333: imageROM = 8'd72;
                4334: imageROM = 8'd37;
                4335: imageROM = 8'd70;
                4336: imageROM = 8'd142;
                4337: imageROM = 8'd73;
                4338: imageROM = 8'd182;
                4339: imageROM = 8'd78;
                4340: imageROM = 8'd30;
                4341: imageROM = 8'd70;
                4342: imageROM = 8'd145;
                4343: imageROM = 8'd73;
                4344: imageROM = 8'd181;
                4345: imageROM = 8'd81;
                4346: imageROM = 8'd26;
                4347: imageROM = 8'd70;
                4348: imageROM = 8'd146;
                4349: imageROM = 8'd74;
                4350: imageROM = 8'd180;
                4351: imageROM = 8'd83;
                4352: imageROM = 8'd23;
                4353: imageROM = 8'd70;
                4354: imageROM = 8'd147;
                4355: imageROM = 8'd77;
                4356: imageROM = 8'd177;
                4357: imageROM = 8'd85;
                4358: imageROM = 8'd20;
                4359: imageROM = 8'd69;
                4360: imageROM = 8'd150;
                4361: imageROM = 8'd81;
                4362: imageROM = 8'd174;
                4363: imageROM = 8'd84;
                4364: imageROM = 8'd18;
                4365: imageROM = 8'd69;
                4366: imageROM = 8'd152;
                4367: imageROM = 8'd79;
                4368: imageROM = 8'd180;
                4369: imageROM = 8'd80;
                4370: imageROM = 8'd16;
                4371: imageROM = 8'd69;
                4372: imageROM = 8'd153;
                4373: imageROM = 8'd78;
                4374: imageROM = 8'd183;
                4375: imageROM = 8'd77;
            // r08.bmp
                4376: imageROM = 8'd63;
                4377: imageROM = 8'd63;
                4378: imageROM = 8'd63;
                4379: imageROM = 8'd63;
                4380: imageROM = 8'd63;
                4381: imageROM = 8'd63;
                4382: imageROM = 8'd63;
                4383: imageROM = 8'd63;
                4384: imageROM = 8'd63;
                4385: imageROM = 8'd63;
                4386: imageROM = 8'd63;
                4387: imageROM = 8'd63;
                4388: imageROM = 8'd63;
                4389: imageROM = 8'd63;
                4390: imageROM = 8'd63;
                4391: imageROM = 8'd63;
                4392: imageROM = 8'd63;
                4393: imageROM = 8'd63;
                4394: imageROM = 8'd63;
                4395: imageROM = 8'd63;
                4396: imageROM = 8'd63;
                4397: imageROM = 8'd63;
                4398: imageROM = 8'd63;
                4399: imageROM = 8'd63;
                4400: imageROM = 8'd63;
                4401: imageROM = 8'd63;
                4402: imageROM = 8'd63;
                4403: imageROM = 8'd63;
                4404: imageROM = 8'd63;
                4405: imageROM = 8'd63;
                4406: imageROM = 8'd63;
                4407: imageROM = 8'd63;
                4408: imageROM = 8'd63;
                4409: imageROM = 8'd63;
                4410: imageROM = 8'd63;
                4411: imageROM = 8'd63;
                4412: imageROM = 8'd63;
                4413: imageROM = 8'd63;
                4414: imageROM = 8'd63;
                4415: imageROM = 8'd63;
                4416: imageROM = 8'd63;
                4417: imageROM = 8'd63;
                4418: imageROM = 8'd63;
                4419: imageROM = 8'd63;
                4420: imageROM = 8'd63;
                4421: imageROM = 8'd47;
                4422: imageROM = 8'd80;
                4423: imageROM = 8'd63;
                4424: imageROM = 8'd44;
                4425: imageROM = 8'd90;
                4426: imageROM = 8'd63;
                4427: imageROM = 8'd36;
                4428: imageROM = 8'd95;
                4429: imageROM = 8'd63;
                4430: imageROM = 8'd32;
                4431: imageROM = 8'd99;
                4432: imageROM = 8'd63;
                4433: imageROM = 8'd29;
                4434: imageROM = 8'd101;
                4435: imageROM = 8'd63;
                4436: imageROM = 8'd26;
                4437: imageROM = 8'd79;
                4438: imageROM = 8'd140;
                4439: imageROM = 8'd78;
                4440: imageROM = 8'd63;
                4441: imageROM = 8'd23;
                4442: imageROM = 8'd74;
                4443: imageROM = 8'd151;
                4444: imageROM = 8'd74;
                4445: imageROM = 8'd63;
                4446: imageROM = 8'd20;
                4447: imageROM = 8'd74;
                4448: imageROM = 8'd156;
                4449: imageROM = 8'd72;
                4450: imageROM = 8'd63;
                4451: imageROM = 8'd18;
                4452: imageROM = 8'd73;
                4453: imageROM = 8'd159;
                4454: imageROM = 8'd71;
                4455: imageROM = 8'd63;
                4456: imageROM = 8'd17;
                4457: imageROM = 8'd72;
                4458: imageROM = 8'd163;
                4459: imageROM = 8'd70;
                4460: imageROM = 8'd63;
                4461: imageROM = 8'd15;
                4462: imageROM = 8'd72;
                4463: imageROM = 8'd164;
                4464: imageROM = 8'd71;
                4465: imageROM = 8'd63;
                4466: imageROM = 8'd13;
                4467: imageROM = 8'd72;
                4468: imageROM = 8'd166;
                4469: imageROM = 8'd70;
                4470: imageROM = 8'd63;
                4471: imageROM = 8'd12;
                4472: imageROM = 8'd71;
                4473: imageROM = 8'd169;
                4474: imageROM = 8'd70;
                4475: imageROM = 8'd63;
                4476: imageROM = 8'd10;
                4477: imageROM = 8'd71;
                4478: imageROM = 8'd171;
                4479: imageROM = 8'd69;
                4480: imageROM = 8'd63;
                4481: imageROM = 8'd9;
                4482: imageROM = 8'd71;
                4483: imageROM = 8'd172;
                4484: imageROM = 8'd70;
                4485: imageROM = 8'd63;
                4486: imageROM = 8'd7;
                4487: imageROM = 8'd71;
                4488: imageROM = 8'd174;
                4489: imageROM = 8'd69;
                4490: imageROM = 8'd63;
                4491: imageROM = 8'd6;
                4492: imageROM = 8'd71;
                4493: imageROM = 8'd175;
                4494: imageROM = 8'd70;
                4495: imageROM = 8'd63;
                4496: imageROM = 8'd4;
                4497: imageROM = 8'd71;
                4498: imageROM = 8'd138;
                4499: imageROM = 8'd68;
                4500: imageROM = 8'd147;
                4501: imageROM = 8'd69;
                4502: imageROM = 8'd138;
                4503: imageROM = 8'd70;
                4504: imageROM = 8'd63;
                4505: imageROM = 8'd3;
                4506: imageROM = 8'd71;
                4507: imageROM = 8'd138;
                4508: imageROM = 8'd70;
                4509: imageROM = 8'd143;
                4510: imageROM = 8'd74;
                4511: imageROM = 8'd135;
                4512: imageROM = 8'd71;
                4513: imageROM = 8'd63;
                4514: imageROM = 8'd2;
                4515: imageROM = 8'd71;
                4516: imageROM = 8'd138;
                4517: imageROM = 8'd72;
                4518: imageROM = 8'd140;
                4519: imageROM = 8'd78;
                4520: imageROM = 8'd132;
                4521: imageROM = 8'd73;
                4522: imageROM = 8'd63;
                4523: imageROM = 8'd71;
                4524: imageROM = 8'd139;
                4525: imageROM = 8'd72;
                4526: imageROM = 8'd139;
                4527: imageROM = 8'd80;
                4528: imageROM = 8'd131;
                4529: imageROM = 8'd73;
                4530: imageROM = 8'd62;
                4531: imageROM = 8'd71;
                4532: imageROM = 8'd140;
                4533: imageROM = 8'd73;
                4534: imageROM = 8'd138;
                4535: imageROM = 8'd81;
                4536: imageROM = 8'd129;
                4537: imageROM = 8'd74;
                4538: imageROM = 8'd62;
                4539: imageROM = 8'd70;
                4540: imageROM = 8'd141;
                4541: imageROM = 8'd73;
                4542: imageROM = 8'd137;
                4543: imageROM = 8'd82;
                4544: imageROM = 8'd130;
                4545: imageROM = 8'd74;
                4546: imageROM = 8'd60;
                4547: imageROM = 8'd71;
                4548: imageROM = 8'd141;
                4549: imageROM = 8'd73;
                4550: imageROM = 8'd136;
                4551: imageROM = 8'd71;
                4552: imageROM = 8'd198;
                4553: imageROM = 8'd82;
                4554: imageROM = 8'd59;
                4555: imageROM = 8'd71;
                4556: imageROM = 8'd142;
                4557: imageROM = 8'd73;
                4558: imageROM = 8'd136;
                4559: imageROM = 8'd70;
                4560: imageROM = 8'd200;
                4561: imageROM = 8'd82;
                4562: imageROM = 8'd57;
                4563: imageROM = 8'd71;
                4564: imageROM = 8'd143;
                4565: imageROM = 8'd73;
                4566: imageROM = 8'd135;
                4567: imageROM = 8'd70;
                4568: imageROM = 8'd202;
                4569: imageROM = 8'd81;
                4570: imageROM = 8'd57;
                4571: imageROM = 8'd70;
                4572: imageROM = 8'd144;
                4573: imageROM = 8'd73;
                4574: imageROM = 8'd135;
                4575: imageROM = 8'd70;
                4576: imageROM = 8'd202;
                4577: imageROM = 8'd82;
                4578: imageROM = 8'd55;
                4579: imageROM = 8'd70;
                4580: imageROM = 8'd146;
                4581: imageROM = 8'd71;
                4582: imageROM = 8'd136;
                4583: imageROM = 8'd70;
                4584: imageROM = 8'd203;
                4585: imageROM = 8'd70;
                4586: imageROM = 8'd130;
                4587: imageROM = 8'd66;
                4588: imageROM = 8'd130;
                4589: imageROM = 8'd69;
                4590: imageROM = 8'd54;
                4591: imageROM = 8'd71;
                4592: imageROM = 8'd147;
                4593: imageROM = 8'd70;
                4594: imageROM = 8'd135;
                4595: imageROM = 8'd70;
                4596: imageROM = 8'd204;
                4597: imageROM = 8'd70;
                4598: imageROM = 8'd134;
                4599: imageROM = 8'd70;
                4600: imageROM = 8'd53;
                4601: imageROM = 8'd70;
                4602: imageROM = 8'd149;
                4603: imageROM = 8'd67;
                4604: imageROM = 8'd137;
                4605: imageROM = 8'd70;
                4606: imageROM = 8'd205;
                4607: imageROM = 8'd69;
                4608: imageROM = 8'd135;
                4609: imageROM = 8'd69;
                4610: imageROM = 8'd52;
                4611: imageROM = 8'd70;
                4612: imageROM = 8'd162;
                4613: imageROM = 8'd70;
                4614: imageROM = 8'd205;
                4615: imageROM = 8'd69;
                4616: imageROM = 8'd135;
                4617: imageROM = 8'd70;
                4618: imageROM = 8'd51;
                4619: imageROM = 8'd69;
                4620: imageROM = 8'd163;
                4621: imageROM = 8'd70;
                4622: imageROM = 8'd205;
                4623: imageROM = 8'd69;
                4624: imageROM = 8'd136;
                4625: imageROM = 8'd69;
                4626: imageROM = 8'd50;
                4627: imageROM = 8'd70;
                4628: imageROM = 8'd163;
                4629: imageROM = 8'd70;
                4630: imageROM = 8'd205;
                4631: imageROM = 8'd70;
                4632: imageROM = 8'd135;
                4633: imageROM = 8'd70;
                4634: imageROM = 8'd49;
                4635: imageROM = 8'd69;
                4636: imageROM = 8'd164;
                4637: imageROM = 8'd70;
                4638: imageROM = 8'd205;
                4639: imageROM = 8'd70;
                4640: imageROM = 8'd135;
                4641: imageROM = 8'd70;
                4642: imageROM = 8'd48;
                4643: imageROM = 8'd70;
                4644: imageROM = 8'd164;
                4645: imageROM = 8'd70;
                4646: imageROM = 8'd205;
                4647: imageROM = 8'd70;
                4648: imageROM = 8'd136;
                4649: imageROM = 8'd70;
                4650: imageROM = 8'd47;
                4651: imageROM = 8'd69;
                4652: imageROM = 8'd165;
                4653: imageROM = 8'd70;
                4654: imageROM = 8'd205;
                4655: imageROM = 8'd70;
                4656: imageROM = 8'd136;
                4657: imageROM = 8'd70;
                4658: imageROM = 8'd46;
                4659: imageROM = 8'd70;
                4660: imageROM = 8'd165;
                4661: imageROM = 8'd70;
                4662: imageROM = 8'd205;
                4663: imageROM = 8'd70;
                4664: imageROM = 8'd137;
                4665: imageROM = 8'd69;
                4666: imageROM = 8'd46;
                4667: imageROM = 8'd69;
                4668: imageROM = 8'd166;
                4669: imageROM = 8'd70;
                4670: imageROM = 8'd205;
                4671: imageROM = 8'd70;
                4672: imageROM = 8'd137;
                4673: imageROM = 8'd70;
                4674: imageROM = 8'd45;
                4675: imageROM = 8'd69;
                4676: imageROM = 8'd166;
                4677: imageROM = 8'd70;
                4678: imageROM = 8'd205;
                4679: imageROM = 8'd70;
                4680: imageROM = 8'd138;
                4681: imageROM = 8'd69;
                4682: imageROM = 8'd44;
                4683: imageROM = 8'd70;
                4684: imageROM = 8'd167;
                4685: imageROM = 8'd69;
                4686: imageROM = 8'd205;
                4687: imageROM = 8'd70;
                4688: imageROM = 8'd138;
                4689: imageROM = 8'd69;
                4690: imageROM = 8'd44;
                4691: imageROM = 8'd70;
                4692: imageROM = 8'd167;
                4693: imageROM = 8'd69;
                4694: imageROM = 8'd205;
                4695: imageROM = 8'd70;
                4696: imageROM = 8'd138;
                4697: imageROM = 8'd69;
                4698: imageROM = 8'd44;
                4699: imageROM = 8'd69;
                4700: imageROM = 8'd168;
                4701: imageROM = 8'd69;
                4702: imageROM = 8'd205;
                4703: imageROM = 8'd70;
                4704: imageROM = 8'd138;
                4705: imageROM = 8'd70;
                4706: imageROM = 8'd43;
                4707: imageROM = 8'd69;
                4708: imageROM = 8'd168;
                4709: imageROM = 8'd70;
                4710: imageROM = 8'd204;
                4711: imageROM = 8'd69;
                4712: imageROM = 8'd140;
                4713: imageROM = 8'd69;
                4714: imageROM = 8'd43;
                4715: imageROM = 8'd69;
                4716: imageROM = 8'd168;
                4717: imageROM = 8'd70;
                4718: imageROM = 8'd204;
                4719: imageROM = 8'd69;
                4720: imageROM = 8'd140;
                4721: imageROM = 8'd69;
                4722: imageROM = 8'd42;
                4723: imageROM = 8'd70;
                4724: imageROM = 8'd169;
                4725: imageROM = 8'd69;
                4726: imageROM = 8'd203;
                4727: imageROM = 8'd70;
                4728: imageROM = 8'd140;
                4729: imageROM = 8'd69;
                4730: imageROM = 8'd42;
                4731: imageROM = 8'd70;
                4732: imageROM = 8'd169;
                4733: imageROM = 8'd69;
                4734: imageROM = 8'd203;
                4735: imageROM = 8'd70;
                4736: imageROM = 8'd140;
                4737: imageROM = 8'd69;
                4738: imageROM = 8'd42;
                4739: imageROM = 8'd70;
                4740: imageROM = 8'd169;
                4741: imageROM = 8'd70;
                4742: imageROM = 8'd202;
                4743: imageROM = 8'd70;
                4744: imageROM = 8'd140;
                4745: imageROM = 8'd69;
                4746: imageROM = 8'd41;
                4747: imageROM = 8'd71;
                4748: imageROM = 8'd169;
                4749: imageROM = 8'd70;
                4750: imageROM = 8'd201;
                4751: imageROM = 8'd70;
                4752: imageROM = 8'd141;
                4753: imageROM = 8'd69;
                4754: imageROM = 8'd41;
                4755: imageROM = 8'd71;
                4756: imageROM = 8'd170;
                4757: imageROM = 8'd70;
                4758: imageROM = 8'd199;
                4759: imageROM = 8'd71;
                4760: imageROM = 8'd141;
                4761: imageROM = 8'd69;
                4762: imageROM = 8'd40;
                4763: imageROM = 8'd72;
                4764: imageROM = 8'd170;
                4765: imageROM = 8'd70;
                4766: imageROM = 8'd199;
                4767: imageROM = 8'd70;
                4768: imageROM = 8'd142;
                4769: imageROM = 8'd69;
                4770: imageROM = 8'd39;
                4771: imageROM = 8'd74;
                4772: imageROM = 8'd170;
                4773: imageROM = 8'd70;
                4774: imageROM = 8'd197;
                4775: imageROM = 8'd71;
                4776: imageROM = 8'd142;
                4777: imageROM = 8'd69;
                4778: imageROM = 8'd38;
                4779: imageROM = 8'd75;
                4780: imageROM = 8'd170;
                4781: imageROM = 8'd71;
                4782: imageROM = 8'd196;
                4783: imageROM = 8'd70;
                4784: imageROM = 8'd143;
                4785: imageROM = 8'd69;
                4786: imageROM = 8'd38;
                4787: imageROM = 8'd75;
                4788: imageROM = 8'd171;
                4789: imageROM = 8'd70;
                4790: imageROM = 8'd195;
                4791: imageROM = 8'd70;
                4792: imageROM = 8'd143;
                4793: imageROM = 8'd69;
                4794: imageROM = 8'd38;
                4795: imageROM = 8'd77;
                4796: imageROM = 8'd171;
                4797: imageROM = 8'd70;
                4798: imageROM = 8'd193;
                4799: imageROM = 8'd71;
                4800: imageROM = 8'd143;
                4801: imageROM = 8'd69;
                4802: imageROM = 8'd37;
                4803: imageROM = 8'd71;
                4804: imageROM = 8'd130;
                4805: imageROM = 8'd69;
                4806: imageROM = 8'd171;
                4807: imageROM = 8'd77;
                4808: imageROM = 8'd143;
                4809: imageROM = 8'd70;
                4810: imageROM = 8'd36;
                4811: imageROM = 8'd71;
                4812: imageROM = 8'd131;
                4813: imageROM = 8'd69;
                4814: imageROM = 8'd172;
                4815: imageROM = 8'd75;
                4816: imageROM = 8'd144;
                4817: imageROM = 8'd69;
                4818: imageROM = 8'd36;
                4819: imageROM = 8'd71;
                4820: imageROM = 8'd132;
                4821: imageROM = 8'd70;
                4822: imageROM = 8'd172;
                4823: imageROM = 8'd74;
                4824: imageROM = 8'd144;
                4825: imageROM = 8'd69;
                4826: imageROM = 8'd35;
                4827: imageROM = 8'd71;
                4828: imageROM = 8'd134;
                4829: imageROM = 8'd69;
                4830: imageROM = 8'd172;
                4831: imageROM = 8'd74;
                4832: imageROM = 8'd143;
                4833: imageROM = 8'd70;
                4834: imageROM = 8'd34;
                4835: imageROM = 8'd71;
                4836: imageROM = 8'd135;
                4837: imageROM = 8'd70;
                4838: imageROM = 8'd172;
                4839: imageROM = 8'd72;
                4840: imageROM = 8'd144;
                4841: imageROM = 8'd70;
                4842: imageROM = 8'd33;
                4843: imageROM = 8'd71;
                4844: imageROM = 8'd137;
                4845: imageROM = 8'd70;
                4846: imageROM = 8'd172;
                4847: imageROM = 8'd70;
                4848: imageROM = 8'd145;
                4849: imageROM = 8'd69;
                4850: imageROM = 8'd33;
                4851: imageROM = 8'd71;
                4852: imageROM = 8'd139;
                4853: imageROM = 8'd70;
                4854: imageROM = 8'd172;
                4855: imageROM = 8'd69;
                4856: imageROM = 8'd145;
                4857: imageROM = 8'd69;
                4858: imageROM = 8'd32;
                4859: imageROM = 8'd71;
                4860: imageROM = 8'd140;
                4861: imageROM = 8'd70;
                4862: imageROM = 8'd172;
                4863: imageROM = 8'd68;
                4864: imageROM = 8'd146;
                4865: imageROM = 8'd69;
                4866: imageROM = 8'd31;
                4867: imageROM = 8'd71;
                4868: imageROM = 8'd142;
                4869: imageROM = 8'd70;
                4870: imageROM = 8'd172;
                4871: imageROM = 8'd67;
                4872: imageROM = 8'd146;
                4873: imageROM = 8'd69;
                4874: imageROM = 8'd30;
                4875: imageROM = 8'd71;
                4876: imageROM = 8'd143;
                4877: imageROM = 8'd71;
                4878: imageROM = 8'd172;
                4879: imageROM = 8'd65;
                4880: imageROM = 8'd147;
                4881: imageROM = 8'd69;
                4882: imageROM = 8'd29;
                4883: imageROM = 8'd71;
                4884: imageROM = 8'd145;
                4885: imageROM = 8'd71;
                4886: imageROM = 8'd191;
                4887: imageROM = 8'd69;
                4888: imageROM = 8'd28;
                4889: imageROM = 8'd71;
                4890: imageROM = 8'd147;
                4891: imageROM = 8'd71;
                4892: imageROM = 8'd190;
                4893: imageROM = 8'd69;
                4894: imageROM = 8'd27;
                4895: imageROM = 8'd71;
                4896: imageROM = 8'd149;
                4897: imageROM = 8'd71;
                4898: imageROM = 8'd189;
                4899: imageROM = 8'd69;
                4900: imageROM = 8'd26;
                4901: imageROM = 8'd71;
                4902: imageROM = 8'd151;
                4903: imageROM = 8'd71;
                4904: imageROM = 8'd188;
                4905: imageROM = 8'd69;
                4906: imageROM = 8'd25;
                4907: imageROM = 8'd71;
                4908: imageROM = 8'd153;
                4909: imageROM = 8'd71;
                4910: imageROM = 8'd187;
                4911: imageROM = 8'd70;
                4912: imageROM = 8'd23;
                4913: imageROM = 8'd71;
                4914: imageROM = 8'd155;
                4915: imageROM = 8'd72;
                4916: imageROM = 8'd185;
                4917: imageROM = 8'd70;
                4918: imageROM = 8'd23;
                4919: imageROM = 8'd70;
                4920: imageROM = 8'd157;
                4921: imageROM = 8'd72;
                4922: imageROM = 8'd185;
                4923: imageROM = 8'd69;
                4924: imageROM = 8'd22;
                4925: imageROM = 8'd71;
                4926: imageROM = 8'd158;
                4927: imageROM = 8'd73;
                4928: imageROM = 8'd183;
                4929: imageROM = 8'd70;
                4930: imageROM = 8'd20;
                4931: imageROM = 8'd71;
                4932: imageROM = 8'd161;
                4933: imageROM = 8'd73;
                4934: imageROM = 8'd182;
                4935: imageROM = 8'd69;
                4936: imageROM = 8'd20;
                4937: imageROM = 8'd70;
                4938: imageROM = 8'd163;
                4939: imageROM = 8'd76;
                4940: imageROM = 8'd178;
                4941: imageROM = 8'd70;
                4942: imageROM = 8'd18;
                4943: imageROM = 8'd71;
                4944: imageROM = 8'd165;
                4945: imageROM = 8'd80;
                4946: imageROM = 8'd173;
                4947: imageROM = 8'd70;
                4948: imageROM = 8'd17;
                4949: imageROM = 8'd70;
                4950: imageROM = 8'd167;
                4951: imageROM = 8'd80;
                4952: imageROM = 8'd172;
                4953: imageROM = 8'd71;
                4954: imageROM = 8'd16;
                4955: imageROM = 8'd69;
                4956: imageROM = 8'd170;
                4957: imageROM = 8'd78;
                4958: imageROM = 8'd173;
                4959: imageROM = 8'd70;
            // r09.bmp
                4960: imageROM = 8'd63;
                4961: imageROM = 8'd63;
                4962: imageROM = 8'd63;
                4963: imageROM = 8'd63;
                4964: imageROM = 8'd63;
                4965: imageROM = 8'd63;
                4966: imageROM = 8'd63;
                4967: imageROM = 8'd63;
                4968: imageROM = 8'd63;
                4969: imageROM = 8'd63;
                4970: imageROM = 8'd63;
                4971: imageROM = 8'd63;
                4972: imageROM = 8'd63;
                4973: imageROM = 8'd63;
                4974: imageROM = 8'd63;
                4975: imageROM = 8'd63;
                4976: imageROM = 8'd63;
                4977: imageROM = 8'd63;
                4978: imageROM = 8'd63;
                4979: imageROM = 8'd63;
                4980: imageROM = 8'd63;
                4981: imageROM = 8'd63;
                4982: imageROM = 8'd63;
                4983: imageROM = 8'd63;
                4984: imageROM = 8'd63;
                4985: imageROM = 8'd63;
                4986: imageROM = 8'd63;
                4987: imageROM = 8'd63;
                4988: imageROM = 8'd63;
                4989: imageROM = 8'd63;
                4990: imageROM = 8'd63;
                4991: imageROM = 8'd63;
                4992: imageROM = 8'd63;
                4993: imageROM = 8'd63;
                4994: imageROM = 8'd63;
                4995: imageROM = 8'd63;
                4996: imageROM = 8'd63;
                4997: imageROM = 8'd63;
                4998: imageROM = 8'd63;
                4999: imageROM = 8'd63;
                5000: imageROM = 8'd63;
                5001: imageROM = 8'd51;
                5002: imageROM = 8'd80;
                5003: imageROM = 8'd63;
                5004: imageROM = 8'd45;
                5005: imageROM = 8'd88;
                5006: imageROM = 8'd63;
                5007: imageROM = 8'd39;
                5008: imageROM = 8'd92;
                5009: imageROM = 8'd63;
                5010: imageROM = 8'd34;
                5011: imageROM = 8'd97;
                5012: imageROM = 8'd63;
                5013: imageROM = 8'd30;
                5014: imageROM = 8'd101;
                5015: imageROM = 8'd63;
                5016: imageROM = 8'd27;
                5017: imageROM = 8'd79;
                5018: imageROM = 8'd138;
                5019: imageROM = 8'd79;
                5020: imageROM = 8'd63;
                5021: imageROM = 8'd23;
                5022: imageROM = 8'd77;
                5023: imageROM = 8'd146;
                5024: imageROM = 8'd76;
                5025: imageROM = 8'd63;
                5026: imageROM = 8'd21;
                5027: imageROM = 8'd75;
                5028: imageROM = 8'd152;
                5029: imageROM = 8'd74;
                5030: imageROM = 8'd63;
                5031: imageROM = 8'd18;
                5032: imageROM = 8'd75;
                5033: imageROM = 8'd156;
                5034: imageROM = 8'd74;
                5035: imageROM = 8'd63;
                5036: imageROM = 8'd15;
                5037: imageROM = 8'd74;
                5038: imageROM = 8'd160;
                5039: imageROM = 8'd73;
                5040: imageROM = 8'd63;
                5041: imageROM = 8'd13;
                5042: imageROM = 8'd73;
                5043: imageROM = 8'd163;
                5044: imageROM = 8'd73;
                5045: imageROM = 8'd63;
                5046: imageROM = 8'd11;
                5047: imageROM = 8'd73;
                5048: imageROM = 8'd166;
                5049: imageROM = 8'd71;
                5050: imageROM = 8'd63;
                5051: imageROM = 8'd9;
                5052: imageROM = 8'd73;
                5053: imageROM = 8'd134;
                5054: imageROM = 8'd68;
                5055: imageROM = 8'd147;
                5056: imageROM = 8'd69;
                5057: imageROM = 8'd135;
                5058: imageROM = 8'd71;
                5059: imageROM = 8'd63;
                5060: imageROM = 8'd7;
                5061: imageROM = 8'd73;
                5062: imageROM = 8'd133;
                5063: imageROM = 8'd71;
                5064: imageROM = 8'd143;
                5065: imageROM = 8'd75;
                5066: imageROM = 8'd133;
                5067: imageROM = 8'd71;
                5068: imageROM = 8'd63;
                5069: imageROM = 8'd5;
                5070: imageROM = 8'd72;
                5071: imageROM = 8'd134;
                5072: imageROM = 8'd73;
                5073: imageROM = 8'd141;
                5074: imageROM = 8'd77;
                5075: imageROM = 8'd132;
                5076: imageROM = 8'd71;
                5077: imageROM = 8'd63;
                5078: imageROM = 8'd4;
                5079: imageROM = 8'd72;
                5080: imageROM = 8'd135;
                5081: imageROM = 8'd73;
                5082: imageROM = 8'd140;
                5083: imageROM = 8'd79;
                5084: imageROM = 8'd130;
                5085: imageROM = 8'd73;
                5086: imageROM = 8'd63;
                5087: imageROM = 8'd2;
                5088: imageROM = 8'd72;
                5089: imageROM = 8'd136;
                5090: imageROM = 8'd74;
                5091: imageROM = 8'd138;
                5092: imageROM = 8'd81;
                5093: imageROM = 8'd129;
                5094: imageROM = 8'd73;
                5095: imageROM = 8'd63;
                5096: imageROM = 8'd1;
                5097: imageROM = 8'd72;
                5098: imageROM = 8'd137;
                5099: imageROM = 8'd74;
                5100: imageROM = 8'd137;
                5101: imageROM = 8'd92;
                5102: imageROM = 8'd63;
                5103: imageROM = 8'd72;
                5104: imageROM = 8'd138;
                5105: imageROM = 8'd74;
                5106: imageROM = 8'd136;
                5107: imageROM = 8'd72;
                5108: imageROM = 8'd197;
                5109: imageROM = 8'd80;
                5110: imageROM = 8'd62;
                5111: imageROM = 8'd72;
                5112: imageROM = 8'd139;
                5113: imageROM = 8'd74;
                5114: imageROM = 8'd136;
                5115: imageROM = 8'd70;
                5116: imageROM = 8'd200;
                5117: imageROM = 8'd80;
                5118: imageROM = 8'd60;
                5119: imageROM = 8'd72;
                5120: imageROM = 8'd140;
                5121: imageROM = 8'd74;
                5122: imageROM = 8'd135;
                5123: imageROM = 8'd71;
                5124: imageROM = 8'd201;
                5125: imageROM = 8'd79;
                5126: imageROM = 8'd59;
                5127: imageROM = 8'd72;
                5128: imageROM = 8'd141;
                5129: imageROM = 8'd74;
                5130: imageROM = 8'd135;
                5131: imageROM = 8'd70;
                5132: imageROM = 8'd203;
                5133: imageROM = 8'd78;
                5134: imageROM = 8'd58;
                5135: imageROM = 8'd72;
                5136: imageROM = 8'd143;
                5137: imageROM = 8'd73;
                5138: imageROM = 8'd135;
                5139: imageROM = 8'd70;
                5140: imageROM = 8'd203;
                5141: imageROM = 8'd78;
                5142: imageROM = 8'd57;
                5143: imageROM = 8'd72;
                5144: imageROM = 8'd145;
                5145: imageROM = 8'd72;
                5146: imageROM = 8'd135;
                5147: imageROM = 8'd69;
                5148: imageROM = 8'd204;
                5149: imageROM = 8'd71;
                5150: imageROM = 8'd129;
                5151: imageROM = 8'd71;
                5152: imageROM = 8'd55;
                5153: imageROM = 8'd72;
                5154: imageROM = 8'd147;
                5155: imageROM = 8'd70;
                5156: imageROM = 8'd135;
                5157: imageROM = 8'd70;
                5158: imageROM = 8'd204;
                5159: imageROM = 8'd70;
                5160: imageROM = 8'd131;
                5161: imageROM = 8'd70;
                5162: imageROM = 8'd54;
                5163: imageROM = 8'd72;
                5164: imageROM = 8'd149;
                5165: imageROM = 8'd68;
                5166: imageROM = 8'd136;
                5167: imageROM = 8'd70;
                5168: imageROM = 8'd205;
                5169: imageROM = 8'd70;
                5170: imageROM = 8'd130;
                5171: imageROM = 8'd70;
                5172: imageROM = 8'd53;
                5173: imageROM = 8'd72;
                5174: imageROM = 8'd162;
                5175: imageROM = 8'd70;
                5176: imageROM = 8'd205;
                5177: imageROM = 8'd70;
                5178: imageROM = 8'd131;
                5179: imageROM = 8'd70;
                5180: imageROM = 8'd52;
                5181: imageROM = 8'd71;
                5182: imageROM = 8'd163;
                5183: imageROM = 8'd70;
                5184: imageROM = 8'd205;
                5185: imageROM = 8'd70;
                5186: imageROM = 8'd131;
                5187: imageROM = 8'd70;
                5188: imageROM = 8'd51;
                5189: imageROM = 8'd71;
                5190: imageROM = 8'd164;
                5191: imageROM = 8'd70;
                5192: imageROM = 8'd206;
                5193: imageROM = 8'd69;
                5194: imageROM = 8'd132;
                5195: imageROM = 8'd70;
                5196: imageROM = 8'd49;
                5197: imageROM = 8'd71;
                5198: imageROM = 8'd165;
                5199: imageROM = 8'd70;
                5200: imageROM = 8'd206;
                5201: imageROM = 8'd69;
                5202: imageROM = 8'd132;
                5203: imageROM = 8'd70;
                5204: imageROM = 8'd48;
                5205: imageROM = 8'd71;
                5206: imageROM = 8'd166;
                5207: imageROM = 8'd70;
                5208: imageROM = 8'd205;
                5209: imageROM = 8'd70;
                5210: imageROM = 8'd132;
                5211: imageROM = 8'd71;
                5212: imageROM = 8'd46;
                5213: imageROM = 8'd72;
                5214: imageROM = 8'd166;
                5215: imageROM = 8'd70;
                5216: imageROM = 8'd206;
                5217: imageROM = 8'd70;
                5218: imageROM = 8'd132;
                5219: imageROM = 8'd70;
                5220: imageROM = 8'd46;
                5221: imageROM = 8'd71;
                5222: imageROM = 8'd167;
                5223: imageROM = 8'd70;
                5224: imageROM = 8'd206;
                5225: imageROM = 8'd70;
                5226: imageROM = 8'd133;
                5227: imageROM = 8'd70;
                5228: imageROM = 8'd44;
                5229: imageROM = 8'd71;
                5230: imageROM = 8'd168;
                5231: imageROM = 8'd70;
                5232: imageROM = 8'd206;
                5233: imageROM = 8'd69;
                5234: imageROM = 8'd134;
                5235: imageROM = 8'd70;
                5236: imageROM = 8'd44;
                5237: imageROM = 8'd70;
                5238: imageROM = 8'd169;
                5239: imageROM = 8'd70;
                5240: imageROM = 8'd205;
                5241: imageROM = 8'd70;
                5242: imageROM = 8'd134;
                5243: imageROM = 8'd70;
                5244: imageROM = 8'd43;
                5245: imageROM = 8'd71;
                5246: imageROM = 8'd169;
                5247: imageROM = 8'd70;
                5248: imageROM = 8'd206;
                5249: imageROM = 8'd69;
                5250: imageROM = 8'd135;
                5251: imageROM = 8'd70;
                5252: imageROM = 8'd41;
                5253: imageROM = 8'd72;
                5254: imageROM = 8'd170;
                5255: imageROM = 8'd69;
                5256: imageROM = 8'd206;
                5257: imageROM = 8'd69;
                5258: imageROM = 8'd135;
                5259: imageROM = 8'd70;
                5260: imageROM = 8'd41;
                5261: imageROM = 8'd72;
                5262: imageROM = 8'd170;
                5263: imageROM = 8'd70;
                5264: imageROM = 8'd204;
                5265: imageROM = 8'd70;
                5266: imageROM = 8'd136;
                5267: imageROM = 8'd70;
                5268: imageROM = 8'd39;
                5269: imageROM = 8'd73;
                5270: imageROM = 8'd170;
                5271: imageROM = 8'd70;
                5272: imageROM = 8'd204;
                5273: imageROM = 8'd70;
                5274: imageROM = 8'd136;
                5275: imageROM = 8'd70;
                5276: imageROM = 8'd39;
                5277: imageROM = 8'd73;
                5278: imageROM = 8'd170;
                5279: imageROM = 8'd70;
                5280: imageROM = 8'd204;
                5281: imageROM = 8'd70;
                5282: imageROM = 8'd137;
                5283: imageROM = 8'd69;
                5284: imageROM = 8'd38;
                5285: imageROM = 8'd74;
                5286: imageROM = 8'd171;
                5287: imageROM = 8'd70;
                5288: imageROM = 8'd202;
                5289: imageROM = 8'd71;
                5290: imageROM = 8'd137;
                5291: imageROM = 8'd70;
                5292: imageROM = 8'd37;
                5293: imageROM = 8'd74;
                5294: imageROM = 8'd171;
                5295: imageROM = 8'd70;
                5296: imageROM = 8'd202;
                5297: imageROM = 8'd70;
                5298: imageROM = 8'd138;
                5299: imageROM = 8'd70;
                5300: imageROM = 8'd36;
                5301: imageROM = 8'd75;
                5302: imageROM = 8'd171;
                5303: imageROM = 8'd70;
                5304: imageROM = 8'd202;
                5305: imageROM = 8'd70;
                5306: imageROM = 8'd138;
                5307: imageROM = 8'd70;
                5308: imageROM = 8'd36;
                5309: imageROM = 8'd75;
                5310: imageROM = 8'd172;
                5311: imageROM = 8'd70;
                5312: imageROM = 8'd200;
                5313: imageROM = 8'd70;
                5314: imageROM = 8'd140;
                5315: imageROM = 8'd69;
                5316: imageROM = 8'd36;
                5317: imageROM = 8'd75;
                5318: imageROM = 8'd172;
                5319: imageROM = 8'd70;
                5320: imageROM = 8'd199;
                5321: imageROM = 8'd71;
                5322: imageROM = 8'd140;
                5323: imageROM = 8'd70;
                5324: imageROM = 8'd34;
                5325: imageROM = 8'd70;
                5326: imageROM = 8'd129;
                5327: imageROM = 8'd69;
                5328: imageROM = 8'd172;
                5329: imageROM = 8'd71;
                5330: imageROM = 8'd198;
                5331: imageROM = 8'd71;
                5332: imageROM = 8'd140;
                5333: imageROM = 8'd70;
                5334: imageROM = 8'd34;
                5335: imageROM = 8'd70;
                5336: imageROM = 8'd129;
                5337: imageROM = 8'd69;
                5338: imageROM = 8'd173;
                5339: imageROM = 8'd71;
                5340: imageROM = 8'd196;
                5341: imageROM = 8'd71;
                5342: imageROM = 8'd141;
                5343: imageROM = 8'd70;
                5344: imageROM = 8'd34;
                5345: imageROM = 8'd69;
                5346: imageROM = 8'd130;
                5347: imageROM = 8'd70;
                5348: imageROM = 8'd172;
                5349: imageROM = 8'd71;
                5350: imageROM = 8'd196;
                5351: imageROM = 8'd70;
                5352: imageROM = 8'd142;
                5353: imageROM = 8'd70;
                5354: imageROM = 8'd34;
                5355: imageROM = 8'd69;
                5356: imageROM = 8'd130;
                5357: imageROM = 8'd70;
                5358: imageROM = 8'd173;
                5359: imageROM = 8'd71;
                5360: imageROM = 8'd194;
                5361: imageROM = 8'd71;
                5362: imageROM = 8'd142;
                5363: imageROM = 8'd70;
                5364: imageROM = 8'd33;
                5365: imageROM = 8'd70;
                5366: imageROM = 8'd131;
                5367: imageROM = 8'd69;
                5368: imageROM = 8'd174;
                5369: imageROM = 8'd71;
                5370: imageROM = 8'd193;
                5371: imageROM = 8'd70;
                5372: imageROM = 8'd143;
                5373: imageROM = 8'd70;
                5374: imageROM = 8'd33;
                5375: imageROM = 8'd70;
                5376: imageROM = 8'd131;
                5377: imageROM = 8'd70;
                5378: imageROM = 8'd174;
                5379: imageROM = 8'd76;
                5380: imageROM = 8'd144;
                5381: imageROM = 8'd70;
                5382: imageROM = 8'd32;
                5383: imageROM = 8'd71;
                5384: imageROM = 8'd131;
                5385: imageROM = 8'd70;
                5386: imageROM = 8'd174;
                5387: imageROM = 8'd76;
                5388: imageROM = 8'd144;
                5389: imageROM = 8'd70;
                5390: imageROM = 8'd32;
                5391: imageROM = 8'd70;
                5392: imageROM = 8'd133;
                5393: imageROM = 8'd70;
                5394: imageROM = 8'd174;
                5395: imageROM = 8'd74;
                5396: imageROM = 8'd145;
                5397: imageROM = 8'd70;
                5398: imageROM = 8'd31;
                5399: imageROM = 8'd71;
                5400: imageROM = 8'd133;
                5401: imageROM = 8'd70;
                5402: imageROM = 8'd175;
                5403: imageROM = 8'd73;
                5404: imageROM = 8'd145;
                5405: imageROM = 8'd70;
                5406: imageROM = 8'd30;
                5407: imageROM = 8'd71;
                5408: imageROM = 8'd135;
                5409: imageROM = 8'd70;
                5410: imageROM = 8'd174;
                5411: imageROM = 8'd72;
                5412: imageROM = 8'd146;
                5413: imageROM = 8'd70;
                5414: imageROM = 8'd30;
                5415: imageROM = 8'd71;
                5416: imageROM = 8'd135;
                5417: imageROM = 8'd70;
                5418: imageROM = 8'd175;
                5419: imageROM = 8'd71;
                5420: imageROM = 8'd146;
                5421: imageROM = 8'd70;
                5422: imageROM = 8'd29;
                5423: imageROM = 8'd71;
                5424: imageROM = 8'd137;
                5425: imageROM = 8'd70;
                5426: imageROM = 8'd175;
                5427: imageROM = 8'd69;
                5428: imageROM = 8'd147;
                5429: imageROM = 8'd69;
                5430: imageROM = 8'd29;
                5431: imageROM = 8'd71;
                5432: imageROM = 8'd138;
                5433: imageROM = 8'd71;
                5434: imageROM = 8'd175;
                5435: imageROM = 8'd68;
                5436: imageROM = 8'd146;
                5437: imageROM = 8'd70;
                5438: imageROM = 8'd28;
                5439: imageROM = 8'd71;
                5440: imageROM = 8'd140;
                5441: imageROM = 8'd70;
                5442: imageROM = 8'd175;
                5443: imageROM = 8'd67;
                5444: imageROM = 8'd147;
                5445: imageROM = 8'd70;
                5446: imageROM = 8'd27;
                5447: imageROM = 8'd71;
                5448: imageROM = 8'd142;
                5449: imageROM = 8'd70;
                5450: imageROM = 8'd175;
                5451: imageROM = 8'd66;
                5452: imageROM = 8'd147;
                5453: imageROM = 8'd70;
                5454: imageROM = 8'd26;
                5455: imageROM = 8'd71;
                5456: imageROM = 8'd143;
                5457: imageROM = 8'd71;
                5458: imageROM = 8'd191;
                5459: imageROM = 8'd131;
                5460: imageROM = 8'd70;
                5461: imageROM = 8'd26;
                5462: imageROM = 8'd71;
                5463: imageROM = 8'd145;
                5464: imageROM = 8'd71;
                5465: imageROM = 8'd191;
                5466: imageROM = 8'd130;
                5467: imageROM = 8'd70;
                5468: imageROM = 8'd25;
                5469: imageROM = 8'd71;
                5470: imageROM = 8'd147;
                5471: imageROM = 8'd71;
                5472: imageROM = 8'd191;
                5473: imageROM = 8'd70;
                5474: imageROM = 8'd24;
                5475: imageROM = 8'd72;
                5476: imageROM = 8'd149;
                5477: imageROM = 8'd71;
                5478: imageROM = 8'd190;
                5479: imageROM = 8'd70;
                5480: imageROM = 8'd23;
                5481: imageROM = 8'd72;
                5482: imageROM = 8'd151;
                5483: imageROM = 8'd72;
                5484: imageROM = 8'd188;
                5485: imageROM = 8'd70;
                5486: imageROM = 8'd22;
                5487: imageROM = 8'd72;
                5488: imageROM = 8'd153;
                5489: imageROM = 8'd72;
                5490: imageROM = 8'd186;
                5491: imageROM = 8'd70;
                5492: imageROM = 8'd22;
                5493: imageROM = 8'd72;
                5494: imageROM = 8'd155;
                5495: imageROM = 8'd73;
                5496: imageROM = 8'd184;
                5497: imageROM = 8'd70;
                5498: imageROM = 8'd21;
                5499: imageROM = 8'd72;
                5500: imageROM = 8'd157;
                5501: imageROM = 8'd74;
                5502: imageROM = 8'd182;
                5503: imageROM = 8'd69;
                5504: imageROM = 8'd21;
                5505: imageROM = 8'd72;
                5506: imageROM = 8'd159;
                5507: imageROM = 8'd76;
                5508: imageROM = 8'd178;
                5509: imageROM = 8'd70;
                5510: imageROM = 8'd20;
                5511: imageROM = 8'd72;
                5512: imageROM = 8'd162;
                5513: imageROM = 8'd81;
                5514: imageROM = 8'd171;
                5515: imageROM = 8'd70;
                5516: imageROM = 8'd19;
                5517: imageROM = 8'd72;
                5518: imageROM = 8'd164;
                5519: imageROM = 8'd80;
                5520: imageROM = 8'd171;
                5521: imageROM = 8'd69;
                5522: imageROM = 8'd19;
                5523: imageROM = 8'd72;
                5524: imageROM = 8'd167;
                5525: imageROM = 8'd78;
                5526: imageROM = 8'd170;
                5527: imageROM = 8'd70;
                5528: imageROM = 8'd18;
                5529: imageROM = 8'd72;
                5530: imageROM = 8'd170;
                5531: imageROM = 8'd76;
                5532: imageROM = 8'd170;
                5533: imageROM = 8'd70;
                5534: imageROM = 8'd17;
                5535: imageROM = 8'd72;
                5536: imageROM = 8'd173;
                5537: imageROM = 8'd74;
                5538: imageROM = 8'd170;
                5539: imageROM = 8'd70;
                5540: imageROM = 8'd16;
                5541: imageROM = 8'd72;
                5542: imageROM = 8'd178;
                5543: imageROM = 8'd70;
                5544: imageROM = 8'd170;
                5545: imageROM = 8'd69;
                5546: imageROM = 8'd17;
                5547: imageROM = 8'd71;
                5548: imageROM = 8'd191;
                5549: imageROM = 8'd164;
                5550: imageROM = 8'd69;
                5551: imageROM = 8'd16;
                5552: imageROM = 8'd71;
                5553: imageROM = 8'd191;
                5554: imageROM = 8'd165;
                5555: imageROM = 8'd69;
                5556: imageROM = 8'd16;
                5557: imageROM = 8'd70;
                5558: imageROM = 8'd191;
                5559: imageROM = 8'd166;
                5560: imageROM = 8'd69;
                5561: imageROM = 8'd15;
                5562: imageROM = 8'd70;
                5563: imageROM = 8'd191;
                5564: imageROM = 8'd167;
                5565: imageROM = 8'd70;
            // r10.bmp
                5566: imageROM = 8'd63;
                5567: imageROM = 8'd63;
                5568: imageROM = 8'd63;
                5569: imageROM = 8'd63;
                5570: imageROM = 8'd63;
                5571: imageROM = 8'd63;
                5572: imageROM = 8'd63;
                5573: imageROM = 8'd63;
                5574: imageROM = 8'd63;
                5575: imageROM = 8'd63;
                5576: imageROM = 8'd63;
                5577: imageROM = 8'd63;
                5578: imageROM = 8'd63;
                5579: imageROM = 8'd63;
                5580: imageROM = 8'd63;
                5581: imageROM = 8'd63;
                5582: imageROM = 8'd63;
                5583: imageROM = 8'd63;
                5584: imageROM = 8'd63;
                5585: imageROM = 8'd63;
                5586: imageROM = 8'd63;
                5587: imageROM = 8'd63;
                5588: imageROM = 8'd63;
                5589: imageROM = 8'd63;
                5590: imageROM = 8'd63;
                5591: imageROM = 8'd42;
                5592: imageROM = 8'd80;
                5593: imageROM = 8'd63;
                5594: imageROM = 8'd44;
                5595: imageROM = 8'd89;
                5596: imageROM = 8'd63;
                5597: imageROM = 8'd38;
                5598: imageROM = 8'd94;
                5599: imageROM = 8'd63;
                5600: imageROM = 8'd32;
                5601: imageROM = 8'd99;
                5602: imageROM = 8'd63;
                5603: imageROM = 8'd29;
                5604: imageROM = 8'd101;
                5605: imageROM = 8'd63;
                5606: imageROM = 8'd26;
                5607: imageROM = 8'd105;
                5608: imageROM = 8'd63;
                5609: imageROM = 8'd22;
                5610: imageROM = 8'd77;
                5611: imageROM = 8'd148;
                5612: imageROM = 8'd75;
                5613: imageROM = 8'd63;
                5614: imageROM = 8'd20;
                5615: imageROM = 8'd75;
                5616: imageROM = 8'd153;
                5617: imageROM = 8'd74;
                5618: imageROM = 8'd63;
                5619: imageROM = 8'd17;
                5620: imageROM = 8'd75;
                5621: imageROM = 8'd157;
                5622: imageROM = 8'd73;
                5623: imageROM = 8'd63;
                5624: imageROM = 8'd15;
                5625: imageROM = 8'd74;
                5626: imageROM = 8'd161;
                5627: imageROM = 8'd72;
                5628: imageROM = 8'd63;
                5629: imageROM = 8'd13;
                5630: imageROM = 8'd73;
                5631: imageROM = 8'd164;
                5632: imageROM = 8'd72;
                5633: imageROM = 8'd63;
                5634: imageROM = 8'd10;
                5635: imageROM = 8'd74;
                5636: imageROM = 8'd166;
                5637: imageROM = 8'd72;
                5638: imageROM = 8'd63;
                5639: imageROM = 8'd8;
                5640: imageROM = 8'd73;
                5641: imageROM = 8'd133;
                5642: imageROM = 8'd70;
                5643: imageROM = 8'd158;
                5644: imageROM = 8'd71;
                5645: imageROM = 8'd63;
                5646: imageROM = 8'd7;
                5647: imageROM = 8'd73;
                5648: imageROM = 8'd132;
                5649: imageROM = 8'd73;
                5650: imageROM = 8'd158;
                5651: imageROM = 8'd71;
                5652: imageROM = 8'd63;
                5653: imageROM = 8'd5;
                5654: imageROM = 8'd73;
                5655: imageROM = 8'd133;
                5656: imageROM = 8'd73;
                5657: imageROM = 8'd148;
                5658: imageROM = 8'd65;
                5659: imageROM = 8'd136;
                5660: imageROM = 8'd73;
                5661: imageROM = 8'd63;
                5662: imageROM = 8'd3;
                5663: imageROM = 8'd72;
                5664: imageROM = 8'd135;
                5665: imageROM = 8'd73;
                5666: imageROM = 8'd142;
                5667: imageROM = 8'd74;
                5668: imageROM = 8'd133;
                5669: imageROM = 8'd73;
                5670: imageROM = 8'd63;
                5671: imageROM = 8'd2;
                5672: imageROM = 8'd72;
                5673: imageROM = 8'd136;
                5674: imageROM = 8'd74;
                5675: imageROM = 8'd140;
                5676: imageROM = 8'd76;
                5677: imageROM = 8'd132;
                5678: imageROM = 8'd74;
                5679: imageROM = 8'd63;
                5680: imageROM = 8'd72;
                5681: imageROM = 8'd137;
                5682: imageROM = 8'd74;
                5683: imageROM = 8'd139;
                5684: imageROM = 8'd78;
                5685: imageROM = 8'd131;
                5686: imageROM = 8'd74;
                5687: imageROM = 8'd62;
                5688: imageROM = 8'd72;
                5689: imageROM = 8'd138;
                5690: imageROM = 8'd74;
                5691: imageROM = 8'd138;
                5692: imageROM = 8'd80;
                5693: imageROM = 8'd130;
                5694: imageROM = 8'd75;
                5695: imageROM = 8'd60;
                5696: imageROM = 8'd72;
                5697: imageROM = 8'd139;
                5698: imageROM = 8'd74;
                5699: imageROM = 8'd137;
                5700: imageROM = 8'd94;
                5701: imageROM = 8'd59;
                5702: imageROM = 8'd72;
                5703: imageROM = 8'd140;
                5704: imageROM = 8'd74;
                5705: imageROM = 8'd136;
                5706: imageROM = 8'd72;
                5707: imageROM = 8'd193;
                5708: imageROM = 8'd66;
                5709: imageROM = 8'd193;
                5710: imageROM = 8'd83;
                5711: imageROM = 8'd58;
                5712: imageROM = 8'd72;
                5713: imageROM = 8'd141;
                5714: imageROM = 8'd74;
                5715: imageROM = 8'd136;
                5716: imageROM = 8'd71;
                5717: imageROM = 8'd198;
                5718: imageROM = 8'd82;
                5719: imageROM = 8'd58;
                5720: imageROM = 8'd71;
                5721: imageROM = 8'd143;
                5722: imageROM = 8'd73;
                5723: imageROM = 8'd135;
                5724: imageROM = 8'd71;
                5725: imageROM = 8'd200;
                5726: imageROM = 8'd71;
                5727: imageROM = 8'd129;
                5728: imageROM = 8'd74;
                5729: imageROM = 8'd56;
                5730: imageROM = 8'd71;
                5731: imageROM = 8'd145;
                5732: imageROM = 8'd71;
                5733: imageROM = 8'd136;
                5734: imageROM = 8'd70;
                5735: imageROM = 8'd202;
                5736: imageROM = 8'd70;
                5737: imageROM = 8'd131;
                5738: imageROM = 8'd65;
                5739: imageROM = 8'd129;
                5740: imageROM = 8'd70;
                5741: imageROM = 8'd55;
                5742: imageROM = 8'd71;
                5743: imageROM = 8'd146;
                5744: imageROM = 8'd71;
                5745: imageROM = 8'd136;
                5746: imageROM = 8'd70;
                5747: imageROM = 8'd203;
                5748: imageROM = 8'd70;
                5749: imageROM = 8'd132;
                5750: imageROM = 8'd70;
                5751: imageROM = 8'd54;
                5752: imageROM = 8'd71;
                5753: imageROM = 8'd161;
                5754: imageROM = 8'd70;
                5755: imageROM = 8'd204;
                5756: imageROM = 8'd70;
                5757: imageROM = 8'd132;
                5758: imageROM = 8'd70;
                5759: imageROM = 8'd53;
                5760: imageROM = 8'd71;
                5761: imageROM = 8'd162;
                5762: imageROM = 8'd70;
                5763: imageROM = 8'd204;
                5764: imageROM = 8'd70;
                5765: imageROM = 8'd132;
                5766: imageROM = 8'd70;
                5767: imageROM = 8'd53;
                5768: imageROM = 8'd71;
                5769: imageROM = 8'd162;
                5770: imageROM = 8'd70;
                5771: imageROM = 8'd205;
                5772: imageROM = 8'd70;
                5773: imageROM = 8'd131;
                5774: imageROM = 8'd70;
                5775: imageROM = 8'd52;
                5776: imageROM = 8'd71;
                5777: imageROM = 8'd163;
                5778: imageROM = 8'd70;
                5779: imageROM = 8'd205;
                5780: imageROM = 8'd70;
                5781: imageROM = 8'd132;
                5782: imageROM = 8'd69;
                5783: imageROM = 8'd51;
                5784: imageROM = 8'd71;
                5785: imageROM = 8'd163;
                5786: imageROM = 8'd71;
                5787: imageROM = 8'd205;
                5788: imageROM = 8'd70;
                5789: imageROM = 8'd132;
                5790: imageROM = 8'd69;
                5791: imageROM = 8'd51;
                5792: imageROM = 8'd70;
                5793: imageROM = 8'd164;
                5794: imageROM = 8'd71;
                5795: imageROM = 8'd205;
                5796: imageROM = 8'd70;
                5797: imageROM = 8'd132;
                5798: imageROM = 8'd70;
                5799: imageROM = 8'd49;
                5800: imageROM = 8'd71;
                5801: imageROM = 8'd164;
                5802: imageROM = 8'd71;
                5803: imageROM = 8'd205;
                5804: imageROM = 8'd71;
                5805: imageROM = 8'd131;
                5806: imageROM = 8'd70;
                5807: imageROM = 8'd48;
                5808: imageROM = 8'd71;
                5809: imageROM = 8'd165;
                5810: imageROM = 8'd71;
                5811: imageROM = 8'd205;
                5812: imageROM = 8'd71;
                5813: imageROM = 8'd132;
                5814: imageROM = 8'd70;
                5815: imageROM = 8'd47;
                5816: imageROM = 8'd70;
                5817: imageROM = 8'd166;
                5818: imageROM = 8'd71;
                5819: imageROM = 8'd205;
                5820: imageROM = 8'd71;
                5821: imageROM = 8'd132;
                5822: imageROM = 8'd70;
                5823: imageROM = 8'd46;
                5824: imageROM = 8'd70;
                5825: imageROM = 8'd167;
                5826: imageROM = 8'd71;
                5827: imageROM = 8'd205;
                5828: imageROM = 8'd71;
                5829: imageROM = 8'd132;
                5830: imageROM = 8'd70;
                5831: imageROM = 8'd45;
                5832: imageROM = 8'd71;
                5833: imageROM = 8'd167;
                5834: imageROM = 8'd71;
                5835: imageROM = 8'd205;
                5836: imageROM = 8'd71;
                5837: imageROM = 8'd133;
                5838: imageROM = 8'd70;
                5839: imageROM = 8'd44;
                5840: imageROM = 8'd70;
                5841: imageROM = 8'd169;
                5842: imageROM = 8'd70;
                5843: imageROM = 8'd205;
                5844: imageROM = 8'd71;
                5845: imageROM = 8'd133;
                5846: imageROM = 8'd70;
                5847: imageROM = 8'd43;
                5848: imageROM = 8'd71;
                5849: imageROM = 8'd169;
                5850: imageROM = 8'd70;
                5851: imageROM = 8'd205;
                5852: imageROM = 8'd71;
                5853: imageROM = 8'd134;
                5854: imageROM = 8'd70;
                5855: imageROM = 8'd42;
                5856: imageROM = 8'd71;
                5857: imageROM = 8'd169;
                5858: imageROM = 8'd70;
                5859: imageROM = 8'd205;
                5860: imageROM = 8'd70;
                5861: imageROM = 8'd135;
                5862: imageROM = 8'd70;
                5863: imageROM = 8'd41;
                5864: imageROM = 8'd71;
                5865: imageROM = 8'd170;
                5866: imageROM = 8'd71;
                5867: imageROM = 8'd204;
                5868: imageROM = 8'd70;
                5869: imageROM = 8'd136;
                5870: imageROM = 8'd70;
                5871: imageROM = 8'd39;
                5872: imageROM = 8'd72;
                5873: imageROM = 8'd171;
                5874: imageROM = 8'd70;
                5875: imageROM = 8'd204;
                5876: imageROM = 8'd70;
                5877: imageROM = 8'd136;
                5878: imageROM = 8'd70;
                5879: imageROM = 8'd39;
                5880: imageROM = 8'd72;
                5881: imageROM = 8'd171;
                5882: imageROM = 8'd70;
                5883: imageROM = 8'd204;
                5884: imageROM = 8'd70;
                5885: imageROM = 8'd137;
                5886: imageROM = 8'd70;
                5887: imageROM = 8'd37;
                5888: imageROM = 8'd73;
                5889: imageROM = 8'd171;
                5890: imageROM = 8'd70;
                5891: imageROM = 8'd203;
                5892: imageROM = 8'd70;
                5893: imageROM = 8'd138;
                5894: imageROM = 8'd70;
                5895: imageROM = 8'd37;
                5896: imageROM = 8'd73;
                5897: imageROM = 8'd172;
                5898: imageROM = 8'd70;
                5899: imageROM = 8'd202;
                5900: imageROM = 8'd70;
                5901: imageROM = 8'd139;
                5902: imageROM = 8'd69;
                5903: imageROM = 8'd36;
                5904: imageROM = 8'd74;
                5905: imageROM = 8'd172;
                5906: imageROM = 8'd70;
                5907: imageROM = 8'd202;
                5908: imageROM = 8'd70;
                5909: imageROM = 8'd139;
                5910: imageROM = 8'd70;
                5911: imageROM = 8'd35;
                5912: imageROM = 8'd74;
                5913: imageROM = 8'd172;
                5914: imageROM = 8'd70;
                5915: imageROM = 8'd201;
                5916: imageROM = 8'd71;
                5917: imageROM = 8'd139;
                5918: imageROM = 8'd70;
                5919: imageROM = 8'd35;
                5920: imageROM = 8'd74;
                5921: imageROM = 8'd173;
                5922: imageROM = 8'd70;
                5923: imageROM = 8'd200;
                5924: imageROM = 8'd70;
                5925: imageROM = 8'd141;
                5926: imageROM = 8'd69;
                5927: imageROM = 8'd34;
                5928: imageROM = 8'd75;
                5929: imageROM = 8'd173;
                5930: imageROM = 8'd71;
                5931: imageROM = 8'd198;
                5932: imageROM = 8'd71;
                5933: imageROM = 8'd141;
                5934: imageROM = 8'd69;
                5935: imageROM = 8'd34;
                5936: imageROM = 8'd76;
                5937: imageROM = 8'd172;
                5938: imageROM = 8'd71;
                5939: imageROM = 8'd197;
                5940: imageROM = 8'd71;
                5941: imageROM = 8'd142;
                5942: imageROM = 8'd70;
                5943: imageROM = 8'd32;
                5944: imageROM = 8'd70;
                5945: imageROM = 8'd129;
                5946: imageROM = 8'd70;
                5947: imageROM = 8'd173;
                5948: imageROM = 8'd71;
                5949: imageROM = 8'd196;
                5950: imageROM = 8'd70;
                5951: imageROM = 8'd143;
                5952: imageROM = 8'd70;
                5953: imageROM = 8'd32;
                5954: imageROM = 8'd70;
                5955: imageROM = 8'd129;
                5956: imageROM = 8'd70;
                5957: imageROM = 8'd174;
                5958: imageROM = 8'd71;
                5959: imageROM = 8'd194;
                5960: imageROM = 8'd71;
                5961: imageROM = 8'd143;
                5962: imageROM = 8'd70;
                5963: imageROM = 8'd32;
                5964: imageROM = 8'd70;
                5965: imageROM = 8'd129;
                5966: imageROM = 8'd70;
                5967: imageROM = 8'd174;
                5968: imageROM = 8'd71;
                5969: imageROM = 8'd194;
                5970: imageROM = 8'd70;
                5971: imageROM = 8'd144;
                5972: imageROM = 8'd70;
                5973: imageROM = 8'd31;
                5974: imageROM = 8'd70;
                5975: imageROM = 8'd131;
                5976: imageROM = 8'd70;
                5977: imageROM = 8'd174;
                5978: imageROM = 8'd78;
                5979: imageROM = 8'd144;
                5980: imageROM = 8'd70;
                5981: imageROM = 8'd31;
                5982: imageROM = 8'd70;
                5983: imageROM = 8'd131;
                5984: imageROM = 8'd70;
                5985: imageROM = 8'd175;
                5986: imageROM = 8'd76;
                5987: imageROM = 8'd145;
                5988: imageROM = 8'd70;
                5989: imageROM = 8'd31;
                5990: imageROM = 8'd70;
                5991: imageROM = 8'd131;
                5992: imageROM = 8'd70;
                5993: imageROM = 8'd176;
                5994: imageROM = 8'd75;
                5995: imageROM = 8'd145;
                5996: imageROM = 8'd70;
                5997: imageROM = 8'd30;
                5998: imageROM = 8'd71;
                5999: imageROM = 8'd132;
                6000: imageROM = 8'd70;
                6001: imageROM = 8'd175;
                6002: imageROM = 8'd74;
                6003: imageROM = 8'd146;
                6004: imageROM = 8'd70;
                6005: imageROM = 8'd30;
                6006: imageROM = 8'd70;
                6007: imageROM = 8'd133;
                6008: imageROM = 8'd70;
                6009: imageROM = 8'd176;
                6010: imageROM = 8'd72;
                6011: imageROM = 8'd147;
                6012: imageROM = 8'd70;
                6013: imageROM = 8'd29;
                6014: imageROM = 8'd71;
                6015: imageROM = 8'd134;
                6016: imageROM = 8'd70;
                6017: imageROM = 8'd176;
                6018: imageROM = 8'd71;
                6019: imageROM = 8'd147;
                6020: imageROM = 8'd69;
                6021: imageROM = 8'd29;
                6022: imageROM = 8'd71;
                6023: imageROM = 8'd135;
                6024: imageROM = 8'd71;
                6025: imageROM = 8'd175;
                6026: imageROM = 8'd70;
                6027: imageROM = 8'd148;
                6028: imageROM = 8'd69;
                6029: imageROM = 8'd29;
                6030: imageROM = 8'd70;
                6031: imageROM = 8'd137;
                6032: imageROM = 8'd70;
                6033: imageROM = 8'd176;
                6034: imageROM = 8'd69;
                6035: imageROM = 8'd147;
                6036: imageROM = 8'd70;
                6037: imageROM = 8'd28;
                6038: imageROM = 8'd71;
                6039: imageROM = 8'd137;
                6040: imageROM = 8'd71;
                6041: imageROM = 8'd176;
                6042: imageROM = 8'd67;
                6043: imageROM = 8'd148;
                6044: imageROM = 8'd70;
                6045: imageROM = 8'd27;
                6046: imageROM = 8'd71;
                6047: imageROM = 8'd139;
                6048: imageROM = 8'd71;
                6049: imageROM = 8'd175;
                6050: imageROM = 8'd67;
                6051: imageROM = 8'd148;
                6052: imageROM = 8'd70;
                6053: imageROM = 8'd26;
                6054: imageROM = 8'd71;
                6055: imageROM = 8'd141;
                6056: imageROM = 8'd70;
                6057: imageROM = 8'd176;
                6058: imageROM = 8'd66;
                6059: imageROM = 8'd147;
                6060: imageROM = 8'd70;
                6061: imageROM = 8'd26;
                6062: imageROM = 8'd71;
                6063: imageROM = 8'd142;
                6064: imageROM = 8'd71;
                6065: imageROM = 8'd191;
                6066: imageROM = 8'd133;
                6067: imageROM = 8'd70;
                6068: imageROM = 8'd25;
                6069: imageROM = 8'd72;
                6070: imageROM = 8'd143;
                6071: imageROM = 8'd71;
                6072: imageROM = 8'd191;
                6073: imageROM = 8'd131;
                6074: imageROM = 8'd70;
                6075: imageROM = 8'd25;
                6076: imageROM = 8'd72;
                6077: imageROM = 8'd145;
                6078: imageROM = 8'd71;
                6079: imageROM = 8'd191;
                6080: imageROM = 8'd130;
                6081: imageROM = 8'd70;
                6082: imageROM = 8'd24;
                6083: imageROM = 8'd72;
                6084: imageROM = 8'd147;
                6085: imageROM = 8'd71;
                6086: imageROM = 8'd191;
                6087: imageROM = 8'd71;
                6088: imageROM = 8'd22;
                6089: imageROM = 8'd73;
                6090: imageROM = 8'd149;
                6091: imageROM = 8'd72;
                6092: imageROM = 8'd189;
                6093: imageROM = 8'd70;
                6094: imageROM = 8'd22;
                6095: imageROM = 8'd73;
                6096: imageROM = 8'd151;
                6097: imageROM = 8'd72;
                6098: imageROM = 8'd187;
                6099: imageROM = 8'd71;
                6100: imageROM = 8'd21;
                6101: imageROM = 8'd72;
                6102: imageROM = 8'd153;
                6103: imageROM = 8'd74;
                6104: imageROM = 8'd185;
                6105: imageROM = 8'd70;
                6106: imageROM = 8'd21;
                6107: imageROM = 8'd72;
                6108: imageROM = 8'd156;
                6109: imageROM = 8'd74;
                6110: imageROM = 8'd182;
                6111: imageROM = 8'd71;
                6112: imageROM = 8'd20;
                6113: imageROM = 8'd72;
                6114: imageROM = 8'd158;
                6115: imageROM = 8'd75;
                6116: imageROM = 8'd180;
                6117: imageROM = 8'd70;
                6118: imageROM = 8'd20;
                6119: imageROM = 8'd72;
                6120: imageROM = 8'd160;
                6121: imageROM = 8'd82;
                6122: imageROM = 8'd171;
                6123: imageROM = 8'd71;
                6124: imageROM = 8'd19;
                6125: imageROM = 8'd72;
                6126: imageROM = 8'd163;
                6127: imageROM = 8'd80;
                6128: imageROM = 8'd171;
                6129: imageROM = 8'd70;
                6130: imageROM = 8'd19;
                6131: imageROM = 8'd72;
                6132: imageROM = 8'd166;
                6133: imageROM = 8'd79;
                6134: imageROM = 8'd170;
                6135: imageROM = 8'd70;
                6136: imageROM = 8'd17;
                6137: imageROM = 8'd72;
                6138: imageROM = 8'd169;
                6139: imageROM = 8'd78;
                6140: imageROM = 8'd169;
                6141: imageROM = 8'd70;
                6142: imageROM = 8'd17;
                6143: imageROM = 8'd72;
                6144: imageROM = 8'd173;
                6145: imageROM = 8'd75;
                6146: imageROM = 8'd169;
                6147: imageROM = 8'd70;
                6148: imageROM = 8'd16;
                6149: imageROM = 8'd72;
                6150: imageROM = 8'd177;
                6151: imageROM = 8'd71;
                6152: imageROM = 8'd170;
                6153: imageROM = 8'd70;
                6154: imageROM = 8'd15;
                6155: imageROM = 8'd72;
                6156: imageROM = 8'd191;
                6157: imageROM = 8'd163;
                6158: imageROM = 8'd70;
                6159: imageROM = 8'd15;
                6160: imageROM = 8'd72;
                6161: imageROM = 8'd191;
                6162: imageROM = 8'd164;
                6163: imageROM = 8'd70;
                6164: imageROM = 8'd15;
                6165: imageROM = 8'd71;
                6166: imageROM = 8'd191;
                6167: imageROM = 8'd165;
                6168: imageROM = 8'd70;
                6169: imageROM = 8'd14;
                6170: imageROM = 8'd71;
                6171: imageROM = 8'd191;
                6172: imageROM = 8'd166;
                6173: imageROM = 8'd70;
                6174: imageROM = 8'd13;
                6175: imageROM = 8'd71;
                6176: imageROM = 8'd191;
                6177: imageROM = 8'd166;
                6178: imageROM = 8'd70;
                6179: imageROM = 8'd13;
                6180: imageROM = 8'd71;
                6181: imageROM = 8'd191;
                6182: imageROM = 8'd167;
                6183: imageROM = 8'd70;
                6184: imageROM = 8'd13;
                6185: imageROM = 8'd70;
                6186: imageROM = 8'd191;
                6187: imageROM = 8'd168;
                6188: imageROM = 8'd70;
                6189: imageROM = 8'd12;
                6190: imageROM = 8'd70;
                6191: imageROM = 8'd191;
                6192: imageROM = 8'd168;
                6193: imageROM = 8'd70;
                6194: imageROM = 8'd13;
                6195: imageROM = 8'd70;
                6196: imageROM = 8'd191;
                6197: imageROM = 8'd168;
                6198: imageROM = 8'd70;

                default: imageROM = 8'd0;
            endcase
        end
    endfunction
endmodule
